##
## LEF for PtnCells ;
## created by Innovus v17.11-s080_1 on Mon Jun 21 17:46:16 2021
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO user_proj_example
  CLASS BLOCK ;
  SIZE 158.2400 BY 156.4000 ;
  FOREIGN user_proj_example 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.212 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 92.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.2358 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 97.728 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.492 LAYER met4  ;
    ANTENNAMAXAREACAR 39.542 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 206.868 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.267073 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 155.4800 158.2400 155.6200 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.737 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.524 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.3058 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 8.19811 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 41.1824 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 154.1200 158.2400 154.2600 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 52.1151 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 244.837 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 152.7600 158.2400 152.9000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0745 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 51.3857 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 252.81 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 151.0600 158.2400 151.2000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7384 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.358 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.504 LAYER met2  ;
    ANTENNAMAXAREACAR 73.8377 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 358.317 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 149.7000 158.2400 149.8400 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5941 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.7445 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 65.723 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 323.77 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 148.3400 158.2400 148.4800 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8353 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.9505 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 40.0159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 195.77 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 146.9800 158.2400 147.1200 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.459 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.069 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 66.5952 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 328.131 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 145.2800 158.2400 145.4200 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3605 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 55.8056 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 274.825 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 143.9200 158.2400 144.0600 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4112 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.83 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 50.797 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 250.81 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 142.2200 158.2400 142.3600 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 26.1764 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 128.034 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 140.8600 158.2400 141.0000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 25.7238 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 125.772 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 139.5000 158.2400 139.6400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6032 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.79 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 45.7683 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 225.667 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 137.8000 158.2400 137.9400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7408 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.36 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 32.2729 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 157.986 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 136.4400 158.2400 136.5800 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.861 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 25.2543 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 123.424 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 135.0800 158.2400 135.2200 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1532 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.422 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 26.2693 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 127.695 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 133.3800 158.2400 133.5200 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.623 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 25.7747 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 126.026 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 132.0200 158.2400 132.1600 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6162 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 19.9129 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 95.4808 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 130.6600 158.2400 130.8000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.2558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.168 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 95.7412 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 509.83 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 128.9600 158.2400 129.1000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 35.9339 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 176.822 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 127.6000 158.2400 127.7400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0265 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9065 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 13.2253 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.2242 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 126.2400 158.2400 126.3800 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.4868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.4 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 35.9061 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 192.6 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 124.8800 158.2400 125.0200 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.352 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 114.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.5848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.256 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 38.0139 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 203.006 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 123.1800 158.2400 123.3200 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1882 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.715 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 16.7558 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 80.604 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 121.8200 158.2400 121.9600 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1925 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.75 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.4868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.4 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 44.0313 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 233.802 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 120.4600 158.2400 120.6000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1676 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.612 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 12.4907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 59.2788 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 118.7600 158.2400 118.9000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.426 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 120.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.9008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 29.5238 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 156.335 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 117.4000 158.2400 117.5400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4145 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.7348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 76.9889 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 407.778 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 116.0400 158.2400 116.1800 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.3608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 157.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 5.55576 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 30.0768 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 114.3400 158.2400 114.4800 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3909 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7285 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 12.1598 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 57.6242 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 112.9800 158.2400 113.1200 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4663 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.6768 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.08 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 77.1085 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 401.564 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 111.6200 158.2400 111.7600 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6479 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.9605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.203 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.4258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.408 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 33.7388 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 177.103 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 109.9200 158.2400 110.0600 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1505 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.7198 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 148.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 7.04141 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 38.1212 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 108.5600 158.2400 108.7000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9373 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.4075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.887 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 111.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.7458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 84.448 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 69.8184 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 372.594 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 107.2000 158.2400 107.3400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1904 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.791 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.7958 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 159.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.1708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 40.361 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 214.646 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 105.5000 158.2400 105.6400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4819 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.1305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.8778 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.152 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 30.7202 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 162.085 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 104.1400 158.2400 104.2800 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.3273 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.3575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.252 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 151.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.2928 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 66.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 53.3578 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 284.719 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 102.4400 158.2400 102.5800 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 3.07576 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 15.5677 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 101.0800 158.2400 101.2200 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.2357 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.8995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.069 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 150.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.7938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 84.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 66.3242 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 354.703 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 99.7200 158.2400 99.8600 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.532 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.1048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.904 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 137.248 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 209.712 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 209.11 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 325.173 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 98.0200 158.2400 98.1600 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1917 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.6795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.755 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 111.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.4388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.144 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 44.9735 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 239.758 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 96.6600 158.2400 96.8000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 95.3000 158.2400 95.4400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 93.6000 158.2400 93.7400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 92.2400 158.2400 92.3800 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 90.8800 158.2400 91.0200 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 89.1800 158.2400 89.3200 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 87.8200 158.2400 87.9600 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 86.4600 158.2400 86.6000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 84.7600 158.2400 84.9000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 83.4000 158.2400 83.5400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 82.0400 158.2400 82.1800 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 80.3400 158.2400 80.4800 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 78.9800 158.2400 79.1200 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 77.6200 158.2400 77.7600 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 75.9200 158.2400 76.0600 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 74.5600 158.2400 74.7000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 73.2000 158.2400 73.3400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 71.5000 158.2400 71.6400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 70.1400 158.2400 70.2800 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 68.7800 158.2400 68.9200 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 67.0800 158.2400 67.2200 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 65.7200 158.2400 65.8600 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 64.3600 158.2400 64.5000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 62.6600 158.2400 62.8000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 61.3000 158.2400 61.4400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 59.9400 158.2400 60.0800 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 58.2400 158.2400 58.3800 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 56.8800 158.2400 57.0200 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 55.5200 158.2400 55.6600 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 53.8200 158.2400 53.9600 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 52.4600 158.2400 52.6000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 51.1000 158.2400 51.2400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.7550 49.4000 158.2400 49.5400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0745 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 45.2404 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 223.741 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 48.0400 158.2400 48.1800 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1022 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.9326 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.248 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 46.6800 158.2400 46.8200 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6243 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.8425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.9176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.168 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 45.3200 158.2400 45.4600 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 43.6200 158.2400 43.7600 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.819 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.4408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 77.488 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 42.2600 158.2400 42.4000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.6368 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.958 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 40.9000 158.2400 41.0400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.224 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.894 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 39.2000 158.2400 39.3400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 37.8400 158.2400 37.9800 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3436 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.557 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.1248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.136 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 36.4800 158.2400 36.6200 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.45 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 34.7800 158.2400 34.9200 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.2144 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.846 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 33.4200 158.2400 33.5600 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.623 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 32.0600 158.2400 32.2000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.51 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.324 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 30.3600 158.2400 30.5000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 29.0000 158.2400 29.1400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.5166 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.239 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 27.6400 158.2400 27.7800 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.962 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.584 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 25.9400 158.2400 26.0800 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.1752 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.65 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 24.5800 158.2400 24.7200 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 23.2200 158.2400 23.3600 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.861 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 21.5200 158.2400 21.6600 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.8052 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.8 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 20.1600 158.2400 20.3000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8996 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.154 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 18.8000 158.2400 18.9400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.8664 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.106 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 17.1000 158.2400 17.2400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.2662 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.105 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 15.7400 158.2400 15.8800 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.3257 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.4025 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 14.3800 158.2400 14.5200 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.8024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.786 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 12.6800 158.2400 12.8200 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.9133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.3405 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 11.3200 158.2400 11.4600 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.5952 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.75 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 9.9600 158.2400 10.1000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.6277 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.9125 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 8.2600 158.2400 8.4000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.8643 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.0955 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 6.9000 158.2400 7.0400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.7239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.3935 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 5.5400 158.2400 5.6800 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.0081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.8145 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 3.8400 158.2400 3.9800 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.914 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.344 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 2.4800 158.2400 2.6200 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.1404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.476 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.7550 1.1200 158.2400 1.2600 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 0.7800 0.4850 0.9200 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 1.4600 0.4850 1.6000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 2.1400 0.4850 2.2800 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 3.1600 0.4850 3.3000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 3.8400 0.4850 3.9800 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 4.5200 0.4850 4.6600 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 5.5400 0.4850 5.6800 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 6.2200 0.4850 6.3600 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 7.2400 0.4850 7.3800 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 7.9200 0.4850 8.0600 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 8.6000 0.4850 8.7400 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 9.6200 0.4850 9.7600 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 10.3000 0.4850 10.4400 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 10.9800 0.4850 11.1200 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 12.0000 0.4850 12.1400 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 12.6800 0.4850 12.8200 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 13.7000 0.4850 13.8400 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 14.3800 0.4850 14.5200 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 15.0600 0.4850 15.2000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 16.0800 0.4850 16.2200 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 16.7600 0.4850 16.9000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 17.7800 0.4850 17.9200 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 18.4600 0.4850 18.6000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 19.1400 0.4850 19.2800 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.1600 0.4850 20.3000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.8400 0.4850 20.9800 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 21.5200 0.4850 21.6600 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 22.5400 0.4850 22.6800 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 23.2200 0.4850 23.3600 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 24.2400 0.4850 24.3800 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 24.9200 0.4850 25.0600 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 25.6000 0.4850 25.7400 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 26.6200 0.4850 26.7600 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 27.3000 0.4850 27.4400 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 27.9800 0.4850 28.1200 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 29.0000 0.4850 29.1400 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 29.6800 0.4850 29.8200 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 30.7000 0.4850 30.8400 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 31.3800 0.4850 31.5200 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 32.0600 0.4850 32.2000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 33.0800 0.4850 33.2200 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 33.7600 0.4850 33.9000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 34.7800 0.4850 34.9200 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 35.4600 0.4850 35.6000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 36.1400 0.4850 36.2800 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 37.1600 0.4850 37.3000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 37.8400 0.4850 37.9800 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 38.5200 0.4850 38.6600 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 39.5400 0.4850 39.6800 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 40.2200 0.4850 40.3600 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 41.2400 0.4850 41.3800 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 41.9200 0.4850 42.0600 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 42.6000 0.4850 42.7400 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 43.6200 0.4850 43.7600 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 44.3000 0.4850 44.4400 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 45.3200 0.4850 45.4600 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 46.0000 0.4850 46.1400 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 46.6800 0.4850 46.8200 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 47.7000 0.4850 47.8400 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 48.3800 0.4850 48.5200 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 49.0600 0.4850 49.2000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 50.0800 0.4850 50.2200 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.2817 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.0115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.4078 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 50.0481 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 247.748 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 50.7600 0.4850 50.9000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9612 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.6508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 158.608 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.492 LAYER met3  ;
    ANTENNAMAXAREACAR 62.1672 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 330.67 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.185772 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 51.7800 0.4850 51.9200 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 79.979 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 396.16 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 52.4600 0.4850 52.6000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3058 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.619 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 24.7818 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 130.259 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 53.1400 0.4850 53.2800 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.4851 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 163.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.936 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 8.7196 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 46.202 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 54.1600 0.4850 54.3000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 81.082 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 401.675 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 54.8400 0.4850 54.9800 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6293 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 36.1618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 193.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.3798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 66.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 61.4808 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 325.826 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 55.5200 0.4850 55.6600 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0742 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.8238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.072 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 138.352 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 211.368 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 224.213 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 399.471 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 56.5400 0.4850 56.6800 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.449 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.966 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 34.528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 184.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.6228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 101 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 21.328 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 35.832 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met5  ;
    ANTENNAMAXAREACAR 97.2954 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 187.632 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 57.2200 0.4850 57.3600 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.314 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 42.6812 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 209.493 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 58.2400 0.4850 58.3800 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.091 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.166 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.3008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.616 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 155.248 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 236.712 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 239.744 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 387.106 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 58.9200 0.4850 59.0600 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0749 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.0955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.6808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.768 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 50.8053 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 269.434 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 59.6000 0.4850 59.7400 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3038 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.358 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.363 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 119.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.0118 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 59.2 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 53.5996 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 282.743 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 60.6200 0.4850 60.7600 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3794 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.736 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.1658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.896 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 142.768 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 217.992 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 232.349 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 418.276 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 61.3000 0.4850 61.4400 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0714 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.294 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.3138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.352 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 119.584 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 183.216 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 190.556 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 325.391 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 62.3200 0.4850 62.4600 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.7795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.496 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2954 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 15.3859 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 84.8747 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 63.0000 0.4850 63.1400 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8657 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.3028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 61.4566 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 316.675 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 63.6800 0.4850 63.8200 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.3685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.3518 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.68 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 71.657 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 378.517 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 64.7000 0.4850 64.8400 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1121 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.0548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.096 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 44.4614 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 233.321 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 65.3800 0.4850 65.5200 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4816 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.247 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.35 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 5.88747 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 30.5414 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 66.0600 0.4850 66.2000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1624 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.651 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.177 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.5796 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 18.8707 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 101.438 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 67.0800 0.4850 67.2200 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2059 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.3398 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.616 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 32.1232 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 168.82 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 67.7600 0.4850 67.9000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2339 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.7688 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.904 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 74.756 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 394.574 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 68.7800 0.4850 68.9200 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.882 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.8348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.256 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 50.6719 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 265.685 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 69.4600 0.4850 69.6000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.236 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.901 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.6048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.696 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 36.3988 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 189.099 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 70.1400 0.4850 70.2800 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1358 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.518 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.5388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.344 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 64.9059 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 338.889 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 71.1600 0.4850 71.3000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5968 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.758 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 3.79798 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.0768 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 71.8400 0.4850 71.9800 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1413 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5985 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 26.9257 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 131.192 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 72.8600 0.4850 73.0000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 29.3721 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 143.424 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 73.5400 0.4850 73.6800 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5823 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8035 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 27.6101 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 134.614 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 74.2200 0.4850 74.3600 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1022 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.4888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.744 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 48.5984 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 252.634 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 75.2400 0.4850 75.3800 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.247 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 10.1778 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.499 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 75.9200 0.4850 76.0600 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5968 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.758 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 13.5499 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.8364 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 76.6000 0.4850 76.7400 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0854 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.018 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 117.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 5.09616 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 26.8525 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 77.6200 0.4850 77.7600 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 78.3000 0.4850 78.4400 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 79.3200 0.4850 79.4600 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 80.0000 0.4850 80.1400 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 80.6800 0.4850 80.8200 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 81.7000 0.4850 81.8400 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 82.3800 0.4850 82.5200 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 83.0600 0.4850 83.2000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 84.0800 0.4850 84.2200 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 84.7600 0.4850 84.9000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 85.7800 0.4850 85.9200 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 86.4600 0.4850 86.6000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 87.1400 0.4850 87.2800 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 88.1600 0.4850 88.3000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 88.8400 0.4850 88.9800 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 89.8600 0.4850 90.0000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 90.5400 0.4850 90.6800 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 91.2200 0.4850 91.3600 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 92.2400 0.4850 92.3800 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 92.9200 0.4850 93.0600 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 93.6000 0.4850 93.7400 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 94.6200 0.4850 94.7600 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 95.3000 0.4850 95.4400 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 96.3200 0.4850 96.4600 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 97.0000 0.4850 97.1400 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 97.6800 0.4850 97.8200 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 98.7000 0.4850 98.8400 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 99.3800 0.4850 99.5200 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 100.4000 0.4850 100.5400 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 101.0800 0.4850 101.2200 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 101.7600 0.4850 101.9000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 102.7800 0.4850 102.9200 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 103.4600 0.4850 103.6000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4064 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.806 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 104.1400 0.4850 104.2800 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 105.1600 0.4850 105.3000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.454 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.044 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 105.8400 0.4850 105.9800 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0742 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.631 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 106.8600 0.4850 107.0000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6094 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.821 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 107.5400 0.4850 107.6800 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7727 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7555 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 108.2200 0.4850 108.3600 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4563 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1735 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 109.2400 0.4850 109.3800 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 109.9200 0.4850 110.0600 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 110.6000 0.4850 110.7400 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.819 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.7778 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.952 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 111.6200 0.4850 111.7600 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0629 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.119 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.9368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.8 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 112.3000 0.4850 112.4400 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 113.3200 0.4850 113.4600 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.93 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.424 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 114.0000 0.4850 114.1400 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.5388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.344 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 114.6800 0.4850 114.8200 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6059 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.7505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.2618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.2 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 115.7000 0.4850 115.8400 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.161 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.5588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.784 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 116.3800 0.4850 116.5200 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6765 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.1565 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 117.4000 0.4850 117.5400 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2884 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.216 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 118.0800 0.4850 118.2200 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9776 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.662 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 118.7600 0.4850 118.9000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3664 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.606 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 119.7800 0.4850 119.9200 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.7291 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.3015 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 120.4600 0.4850 120.6000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.091 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.762 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.6938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.504 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 121.1400 0.4850 121.2800 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.7745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.5158 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.888 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 122.1600 0.4850 122.3000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9464 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.506 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 122.8400 0.4850 122.9800 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 123.8600 0.4850 124.0000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8428 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.988 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 124.5400 0.4850 124.6800 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.274 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 125.2200 0.4850 125.3600 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3605 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 126.2400 0.4850 126.3800 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5754 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.598 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.6368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 126.9200 0.4850 127.0600 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6287 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.0628 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.472 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 127.9400 0.4850 128.0800 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9384 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.466 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 128.6200 0.4850 128.7600 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 129.3000 0.4850 129.4400 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0048 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.798 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 130.3200 0.4850 130.4600 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 131.0000 0.4850 131.1400 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2712 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.13 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 131.6800 0.4850 131.8200 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.469 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.6948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.176 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 132.7000 0.4850 132.8400 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.301 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.0208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.248 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 133.3800 0.4850 133.5200 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 134.4000 0.4850 134.5400 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 135.0800 0.4850 135.2200 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3112 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.33 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 135.7600 0.4850 135.9000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 136.7800 0.4850 136.9200 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.7244 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.396 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 137.4600 0.4850 137.6000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.301 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.344 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.4688 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.304 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 138.1400 0.4850 138.2800 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0658 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.0888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.944 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 139.1600 0.4850 139.3000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.6768 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.158 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 139.8400 0.4850 139.9800 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3744 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.646 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 140.8600 0.4850 141.0000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.513 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.9528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.552 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 141.5400 0.4850 141.6800 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 142.2200 0.4850 142.3600 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0233 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.8905 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 143.2400 0.4850 143.3800 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.1997 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.7725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 143.9200 0.4850 144.0600 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.805 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.8548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 79.696 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 144.9400 0.4850 145.0800 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0686 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.9198 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 117.376 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 145.6200 0.4850 145.7600 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7818 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.63 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.9388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.144 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 146.3000 0.4850 146.4400 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0195 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 147.3200 0.4850 147.4600 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8709 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.1935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.3658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.088 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 148.0000 0.4850 148.1400 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.1689 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.6185 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 148.6800 0.4850 148.8200 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.1349 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.4485 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 149.7000 0.4850 149.8400 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 150.3800 0.4850 150.5200 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3605 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 151.4000 0.4850 151.5400 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 152.0800 0.4850 152.2200 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.3085 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.3165 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 152.7600 0.4850 152.9000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0685 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2345 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.6200 155.9150 0.7600 156.4000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.144 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.6608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.328 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1.0800 155.9150 1.2200 156.4000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.8507 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.0275 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2.0000 155.9150 2.1400 156.4000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3975 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8795 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2.9200 155.9150 3.0600 156.4000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0643 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2135 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 3.8400 155.9150 3.9800 156.4000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5406 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.542 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.4888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.744 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 4.3000 155.9150 4.4400 156.4000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4923 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3535 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 5.2200 155.9150 5.3600 156.4000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.3483 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6335 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 6.1400 155.9150 6.2800 156.4000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.1079 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.4315 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 7.0600 155.9150 7.2000 156.4000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1655 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 7.5200 155.9150 7.6600 156.4000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.1907 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.8455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 8.4400 155.9150 8.5800 156.4000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.9311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.4295 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 9.3600 155.9150 9.5000 156.4000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.7719 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.6335 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 10.2800 155.9150 10.4200 156.4000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.233 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.7648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.216 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 10.7400 155.9150 10.8800 156.4000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1894 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.786 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.1588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.984 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 11.6600 155.9150 11.8000 156.4000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.2689 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.1185 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 12.5800 155.9150 12.7200 156.4000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.0907 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.2275 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 13.5000 155.9150 13.6400 156.4000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.064 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.159 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.738 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.2098 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.256 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 13.9600 155.9150 14.1000 156.4000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.4621 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.0845 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 14.8800 155.9150 15.0200 156.4000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.7075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.3115 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 15.8000 155.9150 15.9400 156.4000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4451 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1175 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 16.7200 155.9150 16.8600 156.4000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8936 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.307 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.5028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.152 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 17.1800 155.9150 17.3200 156.4000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.4271 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.0275 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 18.1000 155.9150 18.2400 156.4000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.462 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.251 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.1598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.656 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 19.0200 155.9150 19.1600 156.4000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4227 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8875 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 19.9400 155.9150 20.0800 156.4000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.6179 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.9815 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 20.4000 155.9150 20.5400 156.4000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.7915 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.8495 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 21.3200 155.9150 21.4600 156.4000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.4215 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.8815 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 22.2400 155.9150 22.3800 156.4000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.6832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.0188 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.904 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 23.1600 155.9150 23.3000 156.4000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3975 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8795 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 23.6200 155.9150 23.7600 156.4000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8519 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0335 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 24.5400 155.9150 24.6800 156.4000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6355 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0695 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 25.4600 155.9150 25.6000 156.4000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.8591 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.1875 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 26.3800 155.9150 26.5200 156.4000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.2983 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.2655 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 27.3000 155.9150 27.4400 156.4000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.7579 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.5635 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 27.7600 155.9150 27.9000 156.4000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.2305 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 115.553 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 43.4923 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 207.277 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 28.6800 155.9150 28.8200 156.4000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7014 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.346 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.407 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 141.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.1786 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 252.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 88.1902 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 460.466 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 29.6000 155.9150 29.7400 156.4000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.6273 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.6745 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 28.5048 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 132.687 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 30.5200 155.9150 30.6600 156.4000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.521 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.444 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.697 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 148.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.3816 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 75.8588 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 398.071 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 30.9800 155.9150 31.1200 156.4000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4495 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.6145 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 16.8659 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.2346 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.65092 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.339 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.608 LAYER met3  ;
    ANTENNAGATEAREA 0.621 LAYER met3  ;
    ANTENNAMAXAREACAR 28.6839 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 137.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.715332 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.0107 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.856 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 42.0851 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 209.112 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 31.9000 155.9150 32.0400 156.4000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.1326 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.223 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.896 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 13.9139 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 69.6089 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.778944 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.4258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.408 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 21.1773 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 108.977 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.778944 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 32.8200 155.9150 32.9600 156.4000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.2785 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 19.4173 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 92.6889 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.2334 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.656 LAYER met3  ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 31.7779 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 160.501 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 33.7400 155.9150 33.8800 156.4000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4662 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.17 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.1946 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 136.52 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.429 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 25.744 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 42.456 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.441 LAYER met5  ;
    ANTENNAMAXAREACAR 58.3764 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 96.2721 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 34.2000 155.9150 34.3400 156.4000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.011 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.894 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.947 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.5994 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 180.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 72.6859 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 369.871 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 35.1200 155.9150 35.2600 156.4000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2882 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.28 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.2147 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 40.0229 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 198.275 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.472349 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 36.0400 155.9150 36.1800 156.4000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.1754 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.264 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met2  ;
    ANTENNAMAXAREACAR 12.568 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 56.404 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.453993 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.328 LAYER met3  ;
    ANTENNAGATEAREA 0.8685 LAYER met3  ;
    ANTENNAMAXAREACAR 14.697 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 68.2958 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.500049 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.2717 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 119.248 LAYER met4  ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 37.0918 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 188.203 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 36.9600 155.9150 37.1000 156.4000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.459 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.134 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.415 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.2668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.56 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 7.0506 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 38.2329 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 37.4200 155.9150 37.5600 156.4000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6694 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.186 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.497 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.0014 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 166.272 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 56.3768 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 291.537 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 38.3400 155.9150 38.4800 156.4000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.137 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.2115 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 178.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 77.7757 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 402.789 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 39.2600 155.9150 39.4000 156.4000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.5731 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 97.4155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.8732 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.256 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met3  ;
    ANTENNAMAXAREACAR 22.9451 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 114.003 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.672786 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.5478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.392 LAYER met4  ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 29.5291 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 149.591 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.672786 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 40.1800 155.9150 40.3200 156.4000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.6814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.01 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 67.8151 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 325.337 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.0075 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.976 LAYER met3  ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 71.8412 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 348.063 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 40.6400 155.9150 40.7800 156.4000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2954 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.316 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.769 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.0034 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 219.616 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 48.6781 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 253.622 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 41.5600 155.9150 41.7000 156.4000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2004 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.841 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.8179 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.824 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met3  ;
    ANTENNAMAXAREACAR 41.3672 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 205.034 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.3488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 151.664 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 79.3174 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 408.065 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 42.4800 155.9150 42.6200 156.4000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5344 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.511 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.909 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.8687 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 138.432 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 32.504 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 166.869 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.381719 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 43.4000 155.9150 43.5400 156.4000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.5 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.5941 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.6144 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 228.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 117.497 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 606.221 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 43.8600 155.9150 44.0000 156.4000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7472 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.7949 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 93.6103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 502.921 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.31746 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.2078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.912 LAYER met4  ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 106.891 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 574.225 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.381719 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 44.7800 155.9150 44.9200 156.4000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.747 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.2035 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 33.0088 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 162.344 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.844157 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 45.7000 155.9150 45.8400 156.4000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.772 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.699 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.402 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.7186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 95.44 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 27.3178 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 138.364 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.592162 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 46.6200 155.9150 46.7600 156.4000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0518 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.8895 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 117.68 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 37.9503 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 190.437 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.536761 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 47.0800 155.9150 47.2200 156.4000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.9541 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 119.417 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met2  ;
    ANTENNAMAXAREACAR 48.681 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 232.974 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 48.0000 155.9150 48.1400 156.4000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4662 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.17 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.1618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 108 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 26.9904 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 144.578 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 48.9200 155.9150 49.0600 156.4000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.878 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.1968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.52 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 15.2808 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 81.9708 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 49.8400 155.9150 49.9800 156.4000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.8435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.6475 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.57 LAYER met2  ;
    ANTENNAMAXAREACAR 29.4999 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 137.281 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 50.3000 155.9150 50.4400 156.4000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.0893 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.8465 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met2  ;
    ANTENNAMAXAREACAR 23.8617 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 108.63 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 51.2200 155.9150 51.3600 156.4000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8722 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.7828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 95.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 23.8056 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 127.593 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 52.1400 155.9150 52.2800 156.4000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2348 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.013 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.3488 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.9017 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 90.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8175 LAYER met4  ;
    ANTENNAMAXAREACAR 44.6981 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 236.949 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 53.0600 155.9150 53.2000 156.4000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.657 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.1736 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 151.2 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1325 LAYER met4  ;
    ANTENNAMAXAREACAR 67.6886 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 339.937 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.1135 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 53.9800 155.9150 54.1200 156.4000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.4400 155.9150 54.5800 156.4000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.3600 155.9150 55.5000 156.4000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.2800 155.9150 56.4200 156.4000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.2000 155.9150 57.3400 156.4000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.6600 155.9150 57.8000 156.4000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.5800 155.9150 58.7200 156.4000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.5000 155.9150 59.6400 156.4000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.4200 155.9150 60.5600 156.4000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.8800 155.9150 61.0200 156.4000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.8000 155.9150 61.9400 156.4000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.7200 155.9150 62.8600 156.4000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.6400 155.9150 63.7800 156.4000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.1000 155.9150 64.2400 156.4000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.0200 155.9150 65.1600 156.4000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.9400 155.9150 66.0800 156.4000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.8600 155.9150 67.0000 156.4000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.3200 155.9150 67.4600 156.4000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.2400 155.9150 68.3800 156.4000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.1600 155.9150 69.3000 156.4000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.0800 155.9150 70.2200 156.4000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.5400 155.9150 70.6800 156.4000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.4600 155.9150 71.6000 156.4000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.3800 155.9150 72.5200 156.4000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.3000 155.9150 73.4400 156.4000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.7600 155.9150 73.9000 156.4000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.6800 155.9150 74.8200 156.4000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.6000 155.9150 75.7400 156.4000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.5200 155.9150 76.6600 156.4000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.9800 155.9150 77.1200 156.4000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.9000 155.9150 78.0400 156.4000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.8200 155.9150 78.9600 156.4000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.7400 155.9150 79.8800 156.4000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.6600 155.9150 80.8000 156.4000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.1200 155.9150 81.2600 156.4000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.0400 155.9150 82.1800 156.4000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.9600 155.9150 83.1000 156.4000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.8800 155.9150 84.0200 156.4000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.3400 155.9150 84.4800 156.4000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.2600 155.9150 85.4000 156.4000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.1800 155.9150 86.3200 156.4000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.1000 155.9150 87.2400 156.4000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.5600 155.9150 87.7000 156.4000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.4800 155.9150 88.6200 156.4000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.4000 155.9150 89.5400 156.4000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.3200 155.9150 90.4600 156.4000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.7800 155.9150 90.9200 156.4000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.7000 155.9150 91.8400 156.4000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.6200 155.9150 92.7600 156.4000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.5400 155.9150 93.6800 156.4000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.0000 155.9150 94.1400 156.4000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.9200 155.9150 95.0600 156.4000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.8400 155.9150 95.9800 156.4000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.7600 155.9150 96.9000 156.4000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.2200 155.9150 97.3600 156.4000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.1400 155.9150 98.2800 156.4000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.0600 155.9150 99.2000 156.4000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.9800 155.9150 100.1200 156.4000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.4400 155.9150 100.5800 156.4000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.3600 155.9150 101.5000 156.4000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.2800 155.9150 102.4200 156.4000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.2000 155.9150 103.3400 156.4000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.6600 155.9150 103.8000 156.4000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3808 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.515 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.6498 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.936 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met4  ;
    ANTENNAMAXAREACAR 72.8748 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 387.491 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.413208 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 104.5800 155.9150 104.7200 156.4000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1795 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.7895 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.315 LAYER met2  ;
    ANTENNAMAXAREACAR 23.1349 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 112.222 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.163175 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 105.5000 155.9150 105.6400 156.4000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5195 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.3715 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 13.8285 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 67.3657 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 106.4200 155.9150 106.5600 156.4000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9737 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.7605 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 12.856 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 62.7414 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 107.3400 155.9150 107.4800 156.4000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.332 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.82283 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.4737 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 107.8000 155.9150 107.9400 156.4000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7599 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.5735 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 16.3659 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 79.598 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 108.7200 155.9150 108.8600 156.4000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9051 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.4175 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 12.4865 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 61.0303 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 109.6400 155.9150 109.7800 156.4000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.977 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.0598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.456 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 13.584 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 71.9172 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 110.5600 155.9150 110.7000 156.4000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4662 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.17 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.2228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 18.0273 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 90.2444 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 111.0200 155.9150 111.1600 156.4000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4475 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.1295 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 17.6226 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 86.7111 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 111.9400 155.9150 112.0800 156.4000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6811 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.2975 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 15.0592 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.7576 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 112.8600 155.9150 113.0000 156.4000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3811 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.7975 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 17.3246 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 85.0848 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 113.7800 155.9150 113.9200 156.4000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3808 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.743 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.4778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 72.352 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 37.9469 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 201.537 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 114.2400 155.9150 114.3800 156.4000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.9211 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.4975 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 16.5592 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.3939 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 115.1600 155.9150 115.3000 156.4000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0307 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.0455 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 14.8612 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 72.7677 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 116.0800 155.9150 116.2200 156.4000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5516 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.597 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.0848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.256 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 15.7998 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 79.0141 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 117.0000 155.9150 117.1400 156.4000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.2562 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.12 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.5908 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.288 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 13.3945 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 70.0222 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 117.4600 155.9150 117.6000 156.4000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.573 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.704 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.0508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.408 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 6.81394 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 34.497 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 118.3800 155.9150 118.5200 156.4000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0477 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.0125 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 12.7745 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 62.2323 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 119.3000 155.9150 119.4400 156.4000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8569 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.0585 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 14.6402 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 71.4242 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 120.2200 155.9150 120.3600 156.4000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1067 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3075 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 4.81293 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.4242 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 120.6800 155.9150 120.8200 156.4000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4551 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.0495 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 13.5976 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 66.3475 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 121.6000 155.9150 121.7400 156.4000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.4535 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 12.9527 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.1232 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 122.5200 155.9150 122.6600 156.4000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2199 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.8735 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 13.1224 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.9717 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 123.4400 155.9150 123.5800 156.4000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6483 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.0155 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 14.0887 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 68.6667 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 123.9000 155.9150 124.0400 156.4000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8695 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.1215 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 14.4347 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 70.5333 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 124.8200 155.9150 124.9600 156.4000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8027 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.7875 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 15.0446 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.4465 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 125.7400 155.9150 125.8800 156.4000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9857 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.7025 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 14.6695 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 71.7071 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 126.6600 155.9150 126.8000 156.4000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.2295 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 13.6135 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 66.2909 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 127.1200 155.9150 127.2600 156.4000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8405 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.9765 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 12.356 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 60.1394 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 128.0400 155.9150 128.1800 156.4000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1907 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.8455 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 22.2939 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 109.931 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 128.9600 155.9150 129.1000 156.4000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.9285 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 12.7406 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 62.0626 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 129.8800 155.9150 130.0200 156.4000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5839 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.6935 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 13.8578 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 67.6485 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 130.3400 155.9150 130.4800 156.4000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4929 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.2385 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 14.1396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 68.9212 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 131.2600 155.9150 131.4000 156.4000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.1800 155.9150 132.3200 156.4000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.1000 155.9150 133.2400 156.4000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.0200 155.9150 134.1600 156.4000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.4800 155.9150 134.6200 156.4000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.4000 155.9150 135.5400 156.4000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.3200 155.9150 136.4600 156.4000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.2400 155.9150 137.3800 156.4000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.7000 155.9150 137.8400 156.4000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.6200 155.9150 138.7600 156.4000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.5400 155.9150 139.6800 156.4000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.4600 155.9150 140.6000 156.4000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.9200 155.9150 141.0600 156.4000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.8400 155.9150 141.9800 156.4000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.7600 155.9150 142.9000 156.4000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.6800 155.9150 143.8200 156.4000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.1400 155.9150 144.2800 156.4000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.0600 155.9150 145.2000 156.4000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.9800 155.9150 146.1200 156.4000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.9000 155.9150 147.0400 156.4000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.3600 155.9150 147.5000 156.4000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.2800 155.9150 148.4200 156.4000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.2000 155.9150 149.3400 156.4000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.1200 155.9150 150.2600 156.4000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.5800 155.9150 150.7200 156.4000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.5000 155.9150 151.6400 156.4000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.4200 155.9150 152.5600 156.4000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.3400 155.9150 153.4800 156.4000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.8000 155.9150 153.9400 156.4000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.7200 155.9150 154.8600 156.4000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.6400 155.9150 155.7800 156.4000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.5600 155.9150 156.7000 156.4000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.0200 155.9150 157.1600 156.4000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.4800 0.0000 157.6200 0.4850 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.1000 0.0000 156.2400 0.4850 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.7200 0.0000 154.8600 0.4850 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.3400 0.0000 153.4800 0.4850 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.9600 0.0000 152.1000 0.4850 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.5800 0.0000 150.7200 0.4850 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.2000 0.0000 149.3400 0.4850 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.8200 0.0000 147.9600 0.4850 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.4400 0.0000 146.5800 0.4850 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.0600 0.0000 145.2000 0.4850 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.6800 0.0000 143.8200 0.4850 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.3000 0.0000 142.4400 0.4850 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.9200 0.0000 141.0600 0.4850 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.5400 0.0000 139.6800 0.4850 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.1600 0.0000 138.3000 0.4850 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.7800 0.0000 136.9200 0.4850 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.4000 0.0000 135.5400 0.4850 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.0200 0.0000 134.1600 0.4850 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.6400 0.0000 132.7800 0.4850 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.2600 0.0000 131.4000 0.4850 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.8800 0.0000 130.0200 0.4850 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.5000 0.0000 128.6400 0.4850 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.1200 0.0000 127.2600 0.4850 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.7400 0.0000 125.8800 0.4850 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.3600 0.0000 124.5000 0.4850 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.9800 0.0000 123.1200 0.4850 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.6000 0.0000 121.7400 0.4850 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.2200 0.0000 120.3600 0.4850 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.8400 0.0000 118.9800 0.4850 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.4600 0.0000 117.6000 0.4850 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.0800 0.0000 116.2200 0.4850 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.7000 0.0000 114.8400 0.4850 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.3200 0.0000 113.4600 0.4850 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.9400 0.0000 112.0800 0.4850 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.5600 0.0000 110.7000 0.4850 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.1800 0.0000 109.3200 0.4850 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.8000 0.0000 107.9400 0.4850 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.4200 0.0000 106.5600 0.4850 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.8123 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.9535 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 105.0400 0.0000 105.1800 0.4850 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.9219 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.5015 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 103.6600 0.0000 103.8000 0.4850 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.0003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.8935 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 102.2800 0.0000 102.4200 0.4850 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.9051 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.4175 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 100.9000 0.0000 101.0400 0.4850 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.1907 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.8455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.5200 0.0000 99.6600 0.4850 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.7287 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.5355 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 98.1400 0.0000 98.2800 0.4850 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.1969 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 115.287 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 37.3541 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 185.647 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 96.7600 0.0000 96.9000 0.4850 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0994 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.299 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.1786 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 252.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 54.3219 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 290.248 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 95.3800 0.0000 95.5200 0.4850 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.5937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.4085 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 16.859 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 83.5455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 94.0000 0.0000 94.1400 0.4850 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.611 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.977 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.3816 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 40.6715 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 217.531 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 92.6200 0.0000 92.7600 0.4850 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6556 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.117 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.0107 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.856 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 13.4012 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 72.0964 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 91.2400 0.0000 91.3800 0.4850 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.1026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.234 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7824 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.4258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.408 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 7.26345 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 39.3681 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 89.8600 0.0000 90.0000 0.4850 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.4439 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.646 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.2334 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.656 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 12.3606 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 67.8126 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 88.4800 0.0000 88.6200 0.4850 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.9951 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.3525 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.441 LAYER met2  ;
    ANTENNAMAXAREACAR 48.6183 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 231.603 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.677211 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.441 LAYER met3  ;
    ANTENNAMAXAREACAR 49.1965 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 235.703 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.767914 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3924 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.776 LAYER met4  ;
    ANTENNAGATEAREA 0.441 LAYER met4  ;
    ANTENNAMAXAREACAR 52.3539 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 244.265 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 2.21916 LAYER via4  ;
    ANTENNADIFFAREA 0.429 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 25.744 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 42.456 LAYER met5  ;
    ANTENNAGATEAREA 0.441 LAYER met5  ;
    ANTENNAMAXAREACAR 110.73 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 340.537 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 87.1000 0.0000 87.2400 0.4850 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.096 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.319 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.9351 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.5994 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 180.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 38.6867 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 207.954 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 85.7200 0.0000 85.8600 0.4850 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.0462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 124.726 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 212.563 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 1048.73 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.2147 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.944 LAYER met3  ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 238.285 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1186.54 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 84.3400 0.0000 84.4800 0.4850 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1132 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.4829 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.2717 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 119.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 22.3949 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 119.907 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 82.9600 0.0000 83.1000 0.4850 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.4537 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7735 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 98.381 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 478.758 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.4078 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.112 LAYER met3  ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 114.991 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 568.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.778944 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.2668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.56 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 122.042 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 606.833 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.778944 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 81.5800 0.0000 81.7200 0.4850 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8756 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.217 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.718 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.0014 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 166.272 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 31.1729 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 167.192 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 80.2000 0.0000 80.3400 0.4850 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2702 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.19 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.2115 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 178.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 44.4598 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 238.372 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 78.3600 0.0000 78.5000 0.4850 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.7595 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 83.9556 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 408.425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.8732 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.256 LAYER met3  ;
    ANTENNAGATEAREA 0.9945 LAYER met3  ;
    ANTENNAMAXAREACAR 98.911 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 489.124 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.765618 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.5478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.392 LAYER met4  ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 105.495 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 524.712 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.765618 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 76.9800 0.0000 77.1200 0.4850 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.7737 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.4915 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 30.0766 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 148.422 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.0075 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.976 LAYER met3  ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 34.1027 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 171.148 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 75.6000 0.0000 75.7400 0.4850 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.0034 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 219.616 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 41.2302 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 220.831 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 74.2200 0.0000 74.3600 0.4850 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.2549 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.8345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.3458 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 75.8151 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 389.222 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.3488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 151.664 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 113.765 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 592.253 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 72.8400 0.0000 72.9800 0.4850 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.5068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.082 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 90.0627 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 437.508 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 106.928 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 531.159 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.8687 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 138.432 LAYER met4  ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 132.94 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 670.356 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 71.4600 0.0000 71.6000 0.4850 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.441 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.044 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.6144 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 228.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 57.0474 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 306.142 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 70.0800 0.0000 70.2200 0.4850 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.1556 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 105.273 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 174.869 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 861.119 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.7949 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.368 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 268.479 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1364.04 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.2078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.912 LAYER met4  ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 281.76 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1435.34 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 68.7000 0.0000 68.8400 0.4850 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.0604 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.033 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 83.3167 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 405.23 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 85.4512 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 419.77 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.2035 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.688 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 104.465 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 522.431 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 67.3200 0.0000 67.4600 0.4850 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.8806 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.016 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 79.8214 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 385.175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 81.8452 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 399.524 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.7186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 95.44 LAYER met4  ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 99.6618 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 495.492 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 65.9400 0.0000 66.0800 0.4850 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.293 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 105.437 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 514.897 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 109.707 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 541.373 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.8895 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 117.68 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 139.01 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 698.91 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 64.5600 0.0000 64.7000 0.4850 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.9205 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 119.151 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met2  ;
    ANTENNAMAXAREACAR 24.0528 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 119.809 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 63.1800 0.0000 63.3200 0.4850 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.1984 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.261 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 36.263 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 170.261 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.640055 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 36.6044 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 172.681 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.693603 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.1618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 108 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 63.5947 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 317.26 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.693603 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 61.8000 0.0000 61.9400 0.4850 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.402 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 76.181 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met2  ;
    ANTENNAMAXAREACAR 24.2642 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 114.757 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.448158 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2641 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAGATEAREA 0.9945 LAYER met3  ;
    ANTENNAMAXAREACAR 24.5297 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 116.599 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.488379 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.1968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.52 LAYER met4  ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 39.8106 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 198.57 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.488379 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 60.4200 0.0000 60.5600 0.4850 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.8099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.3815 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.57 LAYER met2  ;
    ANTENNAMAXAREACAR 22.4735 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 111.196 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 59.0400 0.0000 59.1800 0.4850 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.0557 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.5805 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met2  ;
    ANTENNAMAXAREACAR 12.1224 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 59.91 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 57.6600 0.0000 57.8000 0.4850 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.045 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 74.494 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met2  ;
    ANTENNAMAXAREACAR 31.8795 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 148.343 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.640055 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 32.3226 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 151.331 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.693603 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.7828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 95.312 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 56.1282 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 278.924 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.693603 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 56.2800 0.0000 56.4200 0.4850 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.5564 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 57.267 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 106.082 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 520.627 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.92381 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.8949 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.568 LAYER met3  ;
    ANTENNAGATEAREA 0.57 LAYER met3  ;
    ANTENNAMAXAREACAR 114.669 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 567.237 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.993985 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.9017 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 90.608 LAYER met4  ;
    ANTENNAGATEAREA 0.8175 LAYER met4  ;
    ANTENNAMAXAREACAR 135.344 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 678.073 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.993985 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 54.9000 0.0000 55.0400 0.4850 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0994 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.1736 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 151.2 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1325 LAYER met4  ;
    ANTENNAMAXAREACAR 24.8774 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 133.51 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 53.5200 0.0000 53.6600 0.4850 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.1263 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.5235 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 52.1400 0.0000 52.2800 0.4850 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.3898 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 114.128 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 8.7885 LAYER met2  ;
    ANTENNAMAXAREACAR 2.66141 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 12.9861 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 50.7600 0.0000 50.9000 0.4850 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.3653 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 113.957 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 8.7885 LAYER met2  ;
    ANTENNAMAXAREACAR 15.7518 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 75.9908 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.34404 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 49.3800 0.0000 49.5200 0.4850 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.3457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 113.761 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 8.7885 LAYER met2  ;
    ANTENNAMAXAREACAR 2.65639 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 12.9442 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 48.0000 0.0000 48.1400 0.4850 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8067 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0235 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 46.6200 0.0000 46.7600 0.4850 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 45.2400 0.0000 45.3800 0.4850 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 43.8600 0.0000 44.0000 0.4850 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 42.4800 0.0000 42.6200 0.4850 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 41.1000 0.0000 41.2400 0.4850 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 39.7200 0.0000 39.8600 0.4850 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 38.3400 0.0000 38.4800 0.4850 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 36.9600 0.0000 37.1000 0.4850 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 35.5800 0.0000 35.7200 0.4850 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 34.2000 0.0000 34.3400 0.4850 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 32.8200 0.0000 32.9600 0.4850 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 31.4400 0.0000 31.5800 0.4850 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 30.0600 0.0000 30.2000 0.4850 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 28.6800 0.0000 28.8200 0.4850 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 27.3000 0.0000 27.4400 0.4850 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 25.9200 0.0000 26.0600 0.4850 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 24.5400 0.0000 24.6800 0.4850 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 23.1600 0.0000 23.3000 0.4850 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 21.7800 0.0000 21.9200 0.4850 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 20.4000 0.0000 20.5400 0.4850 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 19.0200 0.0000 19.1600 0.4850 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 17.6400 0.0000 17.7800 0.4850 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 16.2600 0.0000 16.4000 0.4850 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 14.8800 0.0000 15.0200 0.4850 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 13.5000 0.0000 13.6400 0.4850 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 12.1200 0.0000 12.2600 0.4850 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 10.7400 0.0000 10.8800 0.4850 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 9.3600 0.0000 9.5000 0.4850 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 7.9800 0.0000 8.1200 0.4850 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 6.6000 0.0000 6.7400 0.4850 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 5.2200 0.0000 5.3600 0.4850 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 3.8400 0.0000 3.9800 0.4850 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2.4600 0.0000 2.6000 0.4850 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.7969 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.8765 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.6200 0.0000 0.7600 0.4850 ;
    END
  END io_oeb[0]
  PIN irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7915 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 153.7800 0.4850 153.9200 ;
    END
  END irq[2]
  PIN irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0798 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.84 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.2948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.376 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 154.4600 0.4850 154.6000 ;
    END
  END irq[1]
  PIN irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 155.4800 0.4850 155.6200 ;
    END
  END irq[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.0000 39.8800 0.4800 40.3600 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 45.3200 0.4800 45.8000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 50.7600 0.4800 51.2400 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 56.2000 0.4800 56.6800 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 61.6400 0.4800 62.1200 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 67.0800 0.4800 67.5600 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 72.5200 0.4800 73.0000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 77.9600 0.4800 78.4400 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 83.4000 0.4800 83.8800 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 88.8400 0.4800 89.3200 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 94.2800 0.4800 94.7600 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 99.7200 0.4800 100.2000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 105.1600 0.4800 105.6400 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 110.6000 0.4800 111.0800 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 116.0400 0.4800 116.5200 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 39.8800 158.2400 40.3600 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 45.3200 158.2400 45.8000 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 50.7600 158.2400 51.2400 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 56.2000 158.2400 56.6800 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 61.6400 158.2400 62.1200 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 67.0800 158.2400 67.5600 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 72.5200 158.2400 73.0000 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 77.9600 158.2400 78.4400 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 83.4000 158.2400 83.8800 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 88.8400 158.2400 89.3200 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 94.2800 158.2400 94.7600 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 99.7200 158.2400 100.2000 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 105.1600 158.2400 105.6400 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 110.6000 158.2400 111.0800 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 116.0400 158.2400 116.5200 ;
    END
    PORT
      LAYER met4 ;
        RECT 40.0200 0.0000 43.3800 3.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 40.0200 153.0400 43.3800 156.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 67.2200 0.0000 70.5800 3.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 67.2200 153.0400 70.5800 156.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 94.4200 0.0000 97.7800 3.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 94.4200 153.0400 97.7800 156.4000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT 40.0200 0.0000 43.3800 156.4000 ;
        RECT 67.2200 0.0000 70.5800 156.4000 ;
        RECT 94.4200 0.0000 97.7800 156.4000 ;
        RECT 39.8550 77.9600 43.3800 78.4400 ;
        RECT 39.8550 39.8800 43.3800 40.3600 ;
        RECT 39.8550 45.3200 43.3800 45.8000 ;
        RECT 39.8550 50.7600 43.3800 51.2400 ;
        RECT 39.8550 56.2000 43.3800 56.6800 ;
        RECT 39.8550 67.0800 43.3800 67.5600 ;
        RECT 39.8550 72.5200 43.3800 73.0000 ;
        RECT 39.8550 61.6400 43.3800 62.1200 ;
        RECT 39.8550 83.4000 43.3800 83.8800 ;
        RECT 39.8550 88.8400 43.3800 89.3200 ;
        RECT 39.8550 94.2800 43.3800 94.7600 ;
        RECT 39.8550 99.7200 43.3800 100.2000 ;
        RECT 39.8550 110.6000 43.3800 111.0800 ;
        RECT 39.8550 116.0400 43.3800 116.5200 ;
        RECT 39.8550 105.1600 43.3800 105.6400 ;
    END
# end of P/G power stripe data as pin

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.0000 42.6000 0.4800 43.0800 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 48.0400 0.4800 48.5200 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 53.4800 0.4800 53.9600 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 58.9200 0.4800 59.4000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 64.3600 0.4800 64.8400 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 69.8000 0.4800 70.2800 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 75.2400 0.4800 75.7200 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 80.6800 0.4800 81.1600 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 86.1200 0.4800 86.6000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 91.5600 0.4800 92.0400 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 97.0000 0.4800 97.4800 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 102.4400 0.4800 102.9200 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 107.8800 0.4800 108.3600 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 113.3200 0.4800 113.8000 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 42.6000 158.2400 43.0800 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 48.0400 158.2400 48.5200 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 53.4800 158.2400 53.9600 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 58.9200 158.2400 59.4000 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 64.3600 158.2400 64.8400 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 69.8000 158.2400 70.2800 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 75.2400 158.2400 75.7200 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 80.6800 158.2400 81.1600 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 86.1200 158.2400 86.6000 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 91.5600 158.2400 92.0400 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 97.0000 158.2400 97.4800 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 102.4400 158.2400 102.9200 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 107.8800 158.2400 108.3600 ;
    END
    PORT
      LAYER met1 ;
        RECT 157.7600 113.3200 158.2400 113.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.6200 0.0000 56.9800 3.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.6200 153.0400 56.9800 156.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 80.8200 0.0000 84.1800 3.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 80.8200 153.0400 84.1800 156.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.0200 0.0000 111.3800 3.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.0200 153.0400 111.3800 156.4000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT 53.6200 0.0000 56.9800 156.4000 ;
        RECT 80.8200 0.0000 84.1800 156.4000 ;
        RECT 108.0200 0.0000 111.3800 156.4000 ;
    END
# end of P/G power stripe data as pin

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.0000 0.0000 158.2400 156.4000 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 158.2400 156.4000 ;
    LAYER met2 ;
      RECT 0.0000 0.0000 158.2400 156.4000 ;
    LAYER met3 ;
      RECT 0.0000 0.0000 158.2400 156.4000 ;
    LAYER met4 ;
      RECT 0.0000 0.0000 158.2400 156.4000 ;
    LAYER met5 ;
      RECT 0.0000 0.0000 158.2400 156.4000 ;
  END
END user_proj_example

END LIBRARY
