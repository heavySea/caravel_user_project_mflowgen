##
## LEF for PtnCells ;
## created by Innovus v17.11-s080_1 on Thu Jun 10 16:32:49 2021
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO user_proj_example
  CLASS BLOCK ;
  SIZE 150.8800 BY 150.9600 ;
  FOREIGN user_proj_example 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.614 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.3078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.492 LAYER met4  ;
    ANTENNAMAXAREACAR 33.5917 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 174.749 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.267073 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 150.0400 150.8800 150.1800 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 43.5352 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 211.5 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 148.6800 150.8800 148.8200 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.3405 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 49.9933 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 239.651 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 147.3200 150.8800 147.4600 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5108 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.328 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 50.273 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 246.52 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 145.9600 150.8800 146.1000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4768 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.988 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 6.85833 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.2976 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.3268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.88 LAYER met3  ;
    ANTENNAGATEAREA 0.504 LAYER met3  ;
    ANTENNAMAXAREACAR 11.475 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 47.8532 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 144.6000 150.8800 144.7400 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4373 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.9605 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 46.4274 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 224.095 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 143.2400 150.8800 143.3800 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0873 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.2105 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 42.7425 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 206.206 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 141.5400 150.8800 141.6800 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9232 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.39 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 33.8996 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 161.456 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 140.1800 150.8800 140.3200 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3215 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.3815 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 36.6647 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 175.817 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 138.8200 150.8800 138.9600 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3605 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 31.6026 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 155.477 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 137.4600 150.8800 137.6000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 24.6139 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 120.533 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 136.1000 150.8800 136.2400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1494 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.586 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.339 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.7328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 73.712 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 58.7206 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 313.594 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 134.7400 150.8800 134.8800 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7956 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.752 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 4.16141 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.1071 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 133.0400 150.8800 133.1800 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 25.1343 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 123.135 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 131.6800 150.8800 131.8200 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.037 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 16.9978 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 82.1253 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 130.3200 150.8800 130.4600 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 26.3844 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 129.386 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 128.9600 150.8800 129.1000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.4635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.7668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.56 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 60.0034 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 316.471 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 127.6000 150.8800 127.7400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7476 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.459 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 12.5093 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 66.3697 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 125.9000 150.8800 126.0400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0714 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.91 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.9028 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 47.952 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 55.5477 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 294.2 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 124.5400 150.8800 124.6800 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7508 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.41 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 23.8188 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 115.754 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 123.1800 150.8800 123.3200 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2366 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.022 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.169 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 113.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.1578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 30.0988 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 160.564 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 121.8200 150.8800 121.9600 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.563 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.0858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.928 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 41.8657 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 222.147 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 120.4600 150.8800 120.6000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8559 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.229 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.9476 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 35.6188 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 192.202 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 119.1000 150.8800 119.2400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.591 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 120.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.2798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.296 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 35.8184 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 189.388 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 117.4000 150.8800 117.5400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1053 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3005 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.62242 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.7212 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 116.0400 150.8800 116.1800 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1477 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.4358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.3038 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.424 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 35.378 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 189.059 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 114.6800 150.8800 114.8200 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.161 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3924 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.776 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 84.592 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 130.728 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 137.59 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 240.246 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 113.3200 150.8800 113.4600 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0994 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.554 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 126.088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.8158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.488 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 32.6952 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 175.552 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 111.9600 150.8800 112.1000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.951 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.872 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.2668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.56 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 25.8923 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 138.6 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 110.2600 150.8800 110.4000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.912 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.098 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 27.7154 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 134.76 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 108.9000 150.8800 109.0400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.496 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.9826 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.848 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 59.1408 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 317.671 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 107.5400 150.8800 107.6800 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4382 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.03 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.5387 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 142.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 4.86121 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 26.5455 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 106.1800 150.8800 106.3200 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.243 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3924 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.776 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 73.216 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 113.664 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 124.412 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 233.695 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 104.8200 150.8800 104.9600 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.1485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 112.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.3908 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 55.888 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 57.6022 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 307.158 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 103.4600 150.8800 103.6000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3279 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.3605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.7058 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.568 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 33.6851 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 178.154 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 101.7600 150.8800 101.9000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.8138 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3924 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.776 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 46.72 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 73.92 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met5  ;
    ANTENNAMAXAREACAR 234.652 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 524.632 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 100.4000 150.8800 100.5400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.38 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 11.5053 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 54.6626 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 99.0400 150.8800 99.1800 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5576 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.562 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 3.36909 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.4545 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 97.6800 150.8800 97.8200 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7742 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.71 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.413 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 141.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.0358 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 40.9586 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 217.206 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 96.3200 150.8800 96.4600 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2678 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.113 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 2.04343 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.44444 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 94.6200 150.8800 94.7600 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.623 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 80.6455 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 400.392 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 93.2600 150.8800 93.4000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 91.9000 150.8800 92.0400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 90.5400 150.8800 90.6800 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 89.1800 150.8800 89.3200 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 87.8200 150.8800 87.9600 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 86.1200 150.8800 86.2600 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 84.7600 150.8800 84.9000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 83.4000 150.8800 83.5400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 82.0400 150.8800 82.1800 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 80.6800 150.8800 80.8200 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 78.9800 150.8800 79.1200 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 77.6200 150.8800 77.7600 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 76.2600 150.8800 76.4000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 74.9000 150.8800 75.0400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 73.5400 150.8800 73.6800 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 72.1800 150.8800 72.3200 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 70.4800 150.8800 70.6200 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 69.1200 150.8800 69.2600 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 67.7600 150.8800 67.9000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 66.4000 150.8800 66.5400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 65.0400 150.8800 65.1800 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 63.3400 150.8800 63.4800 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 61.9800 150.8800 62.1200 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 60.6200 150.8800 60.7600 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 59.2600 150.8800 59.4000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 57.9000 150.8800 58.0400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 56.5400 150.8800 56.6800 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 54.8400 150.8800 54.9800 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 53.4800 150.8800 53.6200 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 52.1200 150.8800 52.2600 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 50.7600 150.8800 50.9000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 49.4000 150.8800 49.5400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 47.7000 150.8800 47.8400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7963 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.7025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.2928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.032 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 38.9456 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 196.27 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 46.3400 150.8800 46.4800 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 44.9800 150.8800 45.1200 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 43.6200 150.8800 43.7600 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.922 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.384 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 42.2600 150.8800 42.4000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.287 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.274 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.732 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.5608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 62.128 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 40.9000 150.8800 41.0400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.796 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.754 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 39.2000 150.8800 39.3400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.695 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.9268 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.08 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 37.8400 150.8800 37.9800 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 36.4800 150.8800 36.6200 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.1188 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.368 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 35.1200 150.8800 35.2600 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.623 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 33.7600 150.8800 33.9000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.394 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 32.0600 150.8800 32.2000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.794 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.6198 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.776 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 30.7000 150.8800 30.8400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 29.3400 150.8800 29.4800 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 27.9800 150.8800 28.1200 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.346 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.504 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 26.6200 150.8800 26.7600 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.3311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.5475 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 25.2600 150.8800 25.4000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 23.5600 150.8800 23.7000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8904 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.226 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 22.2000 150.8800 22.3400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.0824 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.186 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 20.8400 150.8800 20.9800 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.2168 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.858 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 19.4800 150.8800 19.6200 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.1234 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.391 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 18.1200 150.8800 18.2600 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 16.4200 150.8800 16.5600 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4084 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.816 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 15.0600 150.8800 15.2000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.1668 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.608 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 13.7000 150.8800 13.8400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2481 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0145 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 12.3400 150.8800 12.4800 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.6928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.238 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 10.9800 150.8800 11.1200 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9794 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.553 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 9.6200 150.8800 9.7600 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.8797 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.1725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 7.9200 150.8800 8.0600 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.2952 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.25 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 6.5600 150.8800 6.7000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.3568 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.558 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 5.2000 150.8800 5.3400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.2979 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.2635 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 3.8400 150.8800 3.9800 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6436 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.992 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 2.4800 150.8800 2.6200 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.2612 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.08 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 1.1200 150.8800 1.2600 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 0.7800 0.4850 0.9200 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 1.4600 0.4850 1.6000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 2.1400 0.4850 2.2800 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 2.8200 0.4850 2.9600 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 3.8400 0.4850 3.9800 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 4.5200 0.4850 4.6600 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 5.2000 0.4850 5.3400 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 6.2200 0.4850 6.3600 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 6.9000 0.4850 7.0400 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 7.5800 0.4850 7.7200 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 8.2600 0.4850 8.4000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 9.2800 0.4850 9.4200 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 9.9600 0.4850 10.1000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 10.6400 0.4850 10.7800 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 11.6600 0.4850 11.8000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 12.3400 0.4850 12.4800 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 13.0200 0.4850 13.1600 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 14.0400 0.4850 14.1800 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 14.7200 0.4850 14.8600 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 15.4000 0.4850 15.5400 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 16.0800 0.4850 16.2200 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 17.1000 0.4850 17.2400 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 17.7800 0.4850 17.9200 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 18.4600 0.4850 18.6000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 19.4800 0.4850 19.6200 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.1600 0.4850 20.3000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.8400 0.4850 20.9800 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 21.8600 0.4850 22.0000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 22.5400 0.4850 22.6800 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 23.2200 0.4850 23.3600 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 23.9000 0.4850 24.0400 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 24.9200 0.4850 25.0600 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 25.6000 0.4850 25.7400 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 26.2800 0.4850 26.4200 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 27.3000 0.4850 27.4400 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 27.9800 0.4850 28.1200 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 28.6600 0.4850 28.8000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 29.6800 0.4850 29.8200 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 30.3600 0.4850 30.5000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 31.0400 0.4850 31.1800 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 31.7200 0.4850 31.8600 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 32.7400 0.4850 32.8800 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 33.4200 0.4850 33.5600 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 34.1000 0.4850 34.2400 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 35.1200 0.4850 35.2600 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 35.8000 0.4850 35.9400 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 36.4800 0.4850 36.6200 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 37.5000 0.4850 37.6400 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 38.1800 0.4850 38.3200 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 38.8600 0.4850 39.0000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 39.5400 0.4850 39.6800 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 40.5600 0.4850 40.7000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 41.2400 0.4850 41.3800 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 41.9200 0.4850 42.0600 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 42.9400 0.4850 43.0800 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 43.6200 0.4850 43.7600 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 44.3000 0.4850 44.4400 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 45.3200 0.4850 45.4600 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 46.0000 0.4850 46.1400 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 46.6800 0.4850 46.8200 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 47.3600 0.4850 47.5000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 48.3800 0.4850 48.5200 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.6372 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.842 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 55.6142 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 259.77 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 49.0600 0.4850 49.2000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.916 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.0648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 160.816 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.492 LAYER met3  ;
    ANTENNAMAXAREACAR 63.0418 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 335.186 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.185772 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 49.7400 0.4850 49.8800 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.26 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 13.7228 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 65.4566 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 50.7600 0.4850 50.9000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.6804 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.94 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 32.2408 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 157.093 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 51.4400 0.4850 51.5800 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 69.0933 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 342.487 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 52.1200 0.4850 52.2600 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.5445 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 25.9677 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 126.477 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 52.8000 0.4850 52.9400 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.358 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 36.7838 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 180.285 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 53.8200 0.4850 53.9600 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0175 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.828 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 154.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.8886 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 85.68 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 67.462 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 361.895 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 54.5000 0.4850 54.6400 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8144 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.728 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 28.678 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 139.756 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 55.1800 0.4850 55.3200 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0658 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.135 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.3786 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 98.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 78.5481 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 418.772 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 56.2000 0.4850 56.3400 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9779 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.6105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.2848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.656 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 61.9737 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 328.073 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 56.8800 0.4850 57.0200 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.1905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.2 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 34.3362 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 179.43 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 57.5600 0.4850 57.7000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5654 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.548 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.0328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.52 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 118.48 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 181.56 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 188.81 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 321.477 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 58.5800 0.4850 58.7200 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5783 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.5638 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 115.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.7308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 36.368 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 31.6776 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 169.028 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 59.2600 0.4850 59.4000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0882 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.048 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 125.104 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 191.496 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 198.742 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 338.591 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 59.9400 0.4850 60.0800 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8713 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.3028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 41.8032 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 219.164 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 60.6200 0.4850 60.7600 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3563 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.9996 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.272 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 95.2636 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 502.521 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 61.6400 0.4850 61.7800 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7361 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.4015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.8598 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 54.3713 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 286.586 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 62.3200 0.4850 62.4600 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0809 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.5048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.496 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 58.6881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 310.558 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 63.0000 0.4850 63.1400 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.8578 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 38.8588 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 202.347 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 64.0200 0.4850 64.1600 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0949 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.1078 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 47.3556 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 250.703 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 64.7000 0.4850 64.8400 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.532 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.9828 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 76.4255 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 402.618 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 65.3800 0.4850 65.5200 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 39.0877 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 192.758 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 66.4000 0.4850 66.5400 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.425 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.846 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.391 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 15.7208 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 81.4343 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 67.0800 0.4850 67.2200 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.138 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.411 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.6858 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.128 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 41.0436 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 217.628 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 67.7600 0.4850 67.9000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.776 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.654 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.32 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.8869 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 68.4400 0.4850 68.5800 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 25.6729 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 121.889 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 69.4600 0.4850 69.6000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 25.3741 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 124.313 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 70.1400 0.4850 70.2800 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 27.3853 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 131.343 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 70.8200 0.4850 70.9600 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 27.5873 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 133.246 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 71.8400 0.4850 71.9800 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2595 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.973 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.3398 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.616 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 34.8889 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 183.295 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 72.5200 0.4850 72.6600 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2618 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.148 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.1076 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.848 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 74.1444 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 392.166 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 73.2000 0.4850 73.3400 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1372 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.9598 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.256 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 76.4489 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 405.398 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 74.2200 0.4850 74.3600 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 38.8719 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 190.123 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 74.9000 0.4850 75.0400 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 75.5800 0.4850 75.7200 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 76.2600 0.4850 76.4000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 77.2800 0.4850 77.4200 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 77.9600 0.4850 78.1000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 78.6400 0.4850 78.7800 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 79.6600 0.4850 79.8000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 80.3400 0.4850 80.4800 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 81.0200 0.4850 81.1600 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 82.0400 0.4850 82.1800 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 82.7200 0.4850 82.8600 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 83.4000 0.4850 83.5400 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 84.0800 0.4850 84.2200 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 85.1000 0.4850 85.2400 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 85.7800 0.4850 85.9200 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 86.4600 0.4850 86.6000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 87.4800 0.4850 87.6200 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 88.1600 0.4850 88.3000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 88.8400 0.4850 88.9800 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 89.8600 0.4850 90.0000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 90.5400 0.4850 90.6800 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 91.2200 0.4850 91.3600 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 91.9000 0.4850 92.0400 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 92.9200 0.4850 93.0600 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 93.6000 0.4850 93.7400 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 94.2800 0.4850 94.4200 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 95.3000 0.4850 95.4400 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 95.9800 0.4850 96.1200 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 96.6600 0.4850 96.8000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 97.6800 0.4850 97.8200 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 98.3600 0.4850 98.5000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 99.0400 0.4850 99.1800 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 99.7200 0.4850 99.8600 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.238 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 100.7400 0.4850 100.8800 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0882 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.0158 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.888 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 101.4200 0.4850 101.5600 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.51 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.324 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 102.1000 0.4850 102.2400 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 103.1200 0.4850 103.2600 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 103.8000 0.4850 103.9400 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 104.4800 0.4850 104.6200 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.161 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.6488 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.264 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 105.1600 0.4850 105.3000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.274 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 106.1800 0.4850 106.3200 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0919 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3515 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 106.8600 0.4850 107.0000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 107.5400 0.4850 107.6800 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.3558 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.553 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 108.5600 0.4850 108.7000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 109.2400 0.4850 109.3800 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4388 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.968 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 109.9200 0.4850 110.0600 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 110.9400 0.4850 111.0800 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3605 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 111.6200 0.4850 111.7600 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4148 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.848 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 112.3000 0.4850 112.4400 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0798 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.8008 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.408 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 112.9800 0.4850 113.1200 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 114.0000 0.4850 114.1400 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 114.6800 0.4850 114.8200 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3605 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 115.3600 0.4850 115.5000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6405 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.9235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.3438 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.304 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 116.3800 0.4850 116.5200 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6052 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 117.0600 0.4850 117.2000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5919 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.2378 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.072 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 117.7400 0.4850 117.8800 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 118.7600 0.4850 118.9000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5096 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.269 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 119.4400 0.4850 119.5800 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.498 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 120.1200 0.4850 120.2600 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 120.8000 0.4850 120.9400 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6389 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.5008 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.808 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 121.8200 0.4850 121.9600 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.748 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.514 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 122.5000 0.4850 122.6400 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8501 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.0245 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 123.1800 0.4850 123.3200 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 92.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.5108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.528 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 124.2000 0.4850 124.3400 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.082 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 124.8800 0.4850 125.0200 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9708 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.628 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 125.5600 0.4850 125.7000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3112 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.33 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 126.5800 0.4850 126.7200 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.207 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.8148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.816 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 127.2600 0.4850 127.4000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 127.9400 0.4850 128.0800 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9712 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.63 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 128.6200 0.4850 128.7600 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 129.6400 0.4850 129.7800 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 130.3200 0.4850 130.4600 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1798 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.673 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 131.0000 0.4850 131.1400 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9403 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.4225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.2378 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.072 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 132.0200 0.4850 132.1600 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.619 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.2558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.168 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 132.7000 0.4850 132.8400 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0798 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.096 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.4758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 133.3800 0.4850 133.5200 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9433 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.4375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.7448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.776 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 134.4000 0.4850 134.5400 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.6316 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.932 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 135.0800 0.4850 135.2200 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5492 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.52 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 135.7600 0.4850 135.9000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 136.4400 0.4850 136.5800 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 137.4600 0.4850 137.6000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4632 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.037 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.2268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 138.1400 0.4850 138.2800 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4381 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.9645 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 138.8200 0.4850 138.9600 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.318 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.364 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 139.8400 0.4850 139.9800 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7441 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.8438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.304 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 140.5200 0.4850 140.6600 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3605 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 141.2000 0.4850 141.3400 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3961 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 142.2200 0.4850 142.3600 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3605 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 142.9000 0.4850 143.0400 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 143.5800 0.4850 143.7200 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3605 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 144.2600 0.4850 144.4000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0384 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 145.2800 0.4850 145.4200 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6586 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.185 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 145.9600 0.4850 146.1000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3581 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5645 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 146.6400 0.4850 146.7800 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 147.6600 0.4850 147.8000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0518 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.8276 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.688 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.6200 150.4750 0.7600 150.9600 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4927 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3555 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1.0800 150.4750 1.2200 150.9600 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.31 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.389 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.3876 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2.0000 150.4750 2.1400 150.9600 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.756 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.1838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 54.784 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2.9200 150.4750 3.0600 150.9600 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.6491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.0195 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 3.3800 150.4750 3.5200 150.9600 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.8555 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.0515 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 4.3000 150.4750 4.4400 150.9600 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0518 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.4388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.144 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 5.2200 150.4750 5.3600 150.9600 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.351 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.216 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.2956 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 98.856 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.43675 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 69.904 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 108.696 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 5.6800 150.4750 5.8200 150.9600 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1316 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.497 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.7908 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.688 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 6.6000 150.4750 6.7400 150.9600 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.5819 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.6835 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 7.5200 150.4750 7.6600 150.9600 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1144 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.411 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.5748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.536 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 7.9800 150.4750 8.1200 150.9600 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.0127 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.8375 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 8.9000 150.4750 9.0400 150.9600 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.9007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.2775 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 9.8200 150.4750 9.9600 150.9600 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.692 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.4368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.8 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 10.2800 150.4750 10.4200 150.9600 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8109 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8285 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 11.2000 150.4750 11.3400 150.9600 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.0463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.0055 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 12.1200 150.4750 12.2600 150.9600 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8424 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.986 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 12.5800 150.4750 12.7200 150.9600 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.351 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.6238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78.464 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 13.5000 150.4750 13.6400 150.9600 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7828 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.753 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.129 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.4998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.136 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 14.4200 150.4750 14.5600 150.9600 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.8833 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.0725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 14.8800 150.4750 15.0200 150.9600 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7084 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.381 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.4528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.552 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 15.8000 150.4750 15.9400 150.9600 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.7095 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 16.7200 150.4750 16.8600 150.9600 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6978 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.21 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.5368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 17.1800 150.4750 17.3200 150.9600 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.2783 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.1655 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 18.1000 150.4750 18.2400 150.9600 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.7559 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.5535 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 19.0200 150.4750 19.1600 150.9600 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6058 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.868 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.5268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.28 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 19.4800 150.4750 19.6200 150.9600 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8148 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.913 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.921 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.9528 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 69.552 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 20.4000 150.4750 20.5400 150.9600 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7122 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.8128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.472 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 21.3200 150.4750 21.4600 150.9600 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.3123 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.3355 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 21.7800 150.4750 21.9200 150.9600 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.0603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.0755 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 22.7000 150.4750 22.8400 150.9600 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.43 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.924 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 23.6200 150.4750 23.7600 150.9600 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.5671 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.6095 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 24.0800 150.4750 24.2200 150.9600 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.8027 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.7875 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 25.0000 150.4750 25.1400 150.9600 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.5127 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.4555 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 25.9200 150.4750 26.0600 150.9600 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1206 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.442 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.219 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.4018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 45.28 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 26.3800 150.4750 26.5200 150.9600 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.6228 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.858 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 16.7766 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 74.2527 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 27.3000 150.4750 27.4400 150.9600 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.532 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.263 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.098 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 3.83243 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 22.5586 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 28.2200 150.4750 28.3600 150.9600 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.3074 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 60.914 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 37.4805 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 175.924 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.676598 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 38.0548 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 179.996 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.766688 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.2948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.376 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 67.998 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 340.753 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.766688 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 28.6800 150.4750 28.8200 150.9600 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.842 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.62 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 40.2427 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 189.274 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.676598 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 40.8171 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 193.346 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.766688 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.3778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 61.152 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 66.4427 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 331.076 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.766688 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 29.6000 150.4750 29.7400 150.9600 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.566 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.574 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 32.8739 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 154.039 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 30.5200 150.4750 30.6600 150.9600 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.184 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.749 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.2916 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 64.0342 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 335.345 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 31.4400 150.4750 31.5800 150.9600 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.4796 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 96.775 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 55.6452 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 266.747 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.676598 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.672 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 59.9533 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 290.783 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.676598 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 31.9000 150.4750 32.0400 150.9600 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.5798 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.315 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 28.712 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 137.712 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.287421 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.318 LAYER met3  ;
    ANTENNAMAXAREACAR 29.5009 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 143.398 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.413208 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.2936 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 119.84 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 79.7118 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 413.308 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 32.8200 150.4750 32.9600 150.9600 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5776 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.609 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.677 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.0316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 171.296 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 99.4702 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 518.584 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 33.7400 150.4750 33.8800 150.9600 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.5278 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.898 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 34.8377 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 167.847 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.287421 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAGATEAREA 0.318 LAYER met3  ;
    ANTENNAMAXAREACAR 38.0484 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 186.439 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.413208 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.1468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 59.92 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 63.1538 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 321.394 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.413208 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 34.2000 150.4750 34.3400 150.9600 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2914 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.296 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.4766 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.616 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 60.806 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 307.571 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.678207 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.7166 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.096 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 91.6993 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 474.454 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.678207 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 35.1200 150.4750 35.2600 150.9600 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9722 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.7 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.795 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.04 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.5238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.264 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 21.45 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 115.459 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 36.0400 150.4750 36.1800 150.9600 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0518 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.677 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.8646 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 85.552 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 53.0459 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 278.757 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.413208 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 36.5000 150.4750 36.6400 150.9600 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.2894 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.286 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.8057 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 106.096 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 82.9423 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 438.018 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.413208 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 37.4200 150.4750 37.5600 150.9600 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.351 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.9854 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 140 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 94.665 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 494.595 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 38.3400 150.4750 38.4800 150.9600 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8479 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.9405 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 81.7143 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 396.98 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 83.7381 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 411.329 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.6348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.856 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 105.438 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 528.122 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 38.8000 150.4750 38.9400 150.9600 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8892 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.4411 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.8706 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 197.584 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 88.6699 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 470.276 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.413208 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 39.7200 150.4750 39.8600 150.9600 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.06 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.139 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.702 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.9366 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 85.936 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 70.4276 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 357.792 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.946868 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 40.6400 150.4750 40.7800 150.9600 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.4612 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.942 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 28.0505 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 135.422 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 41.1000 150.4750 41.2400 150.9600 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.6324 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 77.798 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 42.6867 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 203.395 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 42.0200 150.4750 42.1600 150.9600 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.059 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.229 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.9097 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 191.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 111.197 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 589.538 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.413208 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 42.9400 150.4750 43.0800 150.9600 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.1954 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.698 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.6507 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.936 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 24.7349 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 127.42 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.287421 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 43.4000 150.4750 43.5400 150.9600 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.1726 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 110.348 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 66.2502 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 320.873 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.498027 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.7408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.088 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 72.4232 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 354.855 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.498027 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 44.3200 150.4750 44.4600 150.9600 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.4952 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.122 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 33.9164 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 160.252 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 45.2400 150.4750 45.3800 150.9600 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.925 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.464 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.401 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.4945 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 206.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 127.074 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 671.29 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 45.7000 150.4750 45.8400 150.9600 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.694 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 88.214 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 60.1231 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 295.02 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 46.6200 150.4750 46.7600 150.9600 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2074 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.876 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.6824 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 154.384 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 82.6198 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 436.712 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 47.5400 150.4750 47.6800 150.9600 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.243 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 27.2849 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 131.197 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.287421 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAGATEAREA 0.318 LAYER met3  ;
    ANTENNAMAXAREACAR 28.1307 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 136.958 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.413208 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.6568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 30.64 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 40.8712 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 205.967 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.413208 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 48.0000 150.4750 48.1400 150.9600 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.5414 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 92.225 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 50.2988 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 240.333 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 48.9200 150.4750 49.0600 150.9600 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.351 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.2968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 108.72 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 45.7135 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 244.865 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 49.8400 150.4750 49.9800 150.9600 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.994 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.724 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 33.4699 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 157.577 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 50.3000 150.4750 50.4400 150.9600 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4732 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.471 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.4633 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 206.544 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.109 LAYER met4  ;
    ANTENNAMAXAREACAR 42.89 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 221.279 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 51.2200 150.4750 51.3600 150.9600 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.1400 150.4750 52.2800 150.9600 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.6000 150.4750 52.7400 150.9600 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.5200 150.4750 53.6600 150.9600 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.4400 150.4750 54.5800 150.9600 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.9000 150.4750 55.0400 150.9600 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.8200 150.4750 55.9600 150.9600 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.7400 150.4750 56.8800 150.9600 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.2000 150.4750 57.3400 150.9600 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.1200 150.4750 58.2600 150.9600 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.0400 150.4750 59.1800 150.9600 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.5000 150.4750 59.6400 150.9600 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.4200 150.4750 60.5600 150.9600 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.3400 150.4750 61.4800 150.9600 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.2600 150.4750 62.4000 150.9600 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.7200 150.4750 62.8600 150.9600 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.6400 150.4750 63.7800 150.9600 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.5600 150.4750 64.7000 150.9600 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.0200 150.4750 65.1600 150.9600 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.9400 150.4750 66.0800 150.9600 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.8600 150.4750 67.0000 150.9600 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.3200 150.4750 67.4600 150.9600 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.2400 150.4750 68.3800 150.9600 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.1600 150.4750 69.3000 150.9600 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.6200 150.4750 69.7600 150.9600 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.5400 150.4750 70.6800 150.9600 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.4600 150.4750 71.6000 150.9600 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.9200 150.4750 72.0600 150.9600 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.8400 150.4750 72.9800 150.9600 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.7600 150.4750 73.9000 150.9600 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.2200 150.4750 74.3600 150.9600 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.1400 150.4750 75.2800 150.9600 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.0600 150.4750 76.2000 150.9600 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.5200 150.4750 76.6600 150.9600 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.4400 150.4750 77.5800 150.9600 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.3600 150.4750 78.5000 150.9600 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.8200 150.4750 78.9600 150.9600 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.7400 150.4750 79.8800 150.9600 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.6600 150.4750 80.8000 150.9600 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.1200 150.4750 81.2600 150.9600 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.0400 150.4750 82.1800 150.9600 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.9600 150.4750 83.1000 150.9600 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.4200 150.4750 83.5600 150.9600 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.3400 150.4750 84.4800 150.9600 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.2600 150.4750 85.4000 150.9600 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.7200 150.4750 85.8600 150.9600 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.6400 150.4750 86.7800 150.9600 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.5600 150.4750 87.7000 150.9600 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.0200 150.4750 88.1600 150.9600 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.9400 150.4750 89.0800 150.9600 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.8600 150.4750 90.0000 150.9600 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.7800 150.4750 90.9200 150.9600 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.2400 150.4750 91.3800 150.9600 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.1600 150.4750 92.3000 150.9600 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.0800 150.4750 93.2200 150.9600 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.5400 150.4750 93.6800 150.9600 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.4600 150.4750 94.6000 150.9600 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.3800 150.4750 95.5200 150.9600 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.8400 150.4750 95.9800 150.9600 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.7600 150.4750 96.9000 150.9600 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.6800 150.4750 97.8200 150.9600 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.1400 150.4750 98.2800 150.9600 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.0600 150.4750 99.2000 150.9600 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3878 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.778 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.7978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 111.392 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met4  ;
    ANTENNAMAXAREACAR 71.0101 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 377.648 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.413208 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 99.9800 150.4750 100.1200 150.9600 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.071 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.194 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.043 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.4888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 61.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.665 LAYER met4  ;
    ANTENNAMAXAREACAR 20.4168 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 107.332 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.197594 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 100.4400 150.4750 100.5800 150.9600 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.2187 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.8675 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 39.5273 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 195.127 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 101.3600 150.4750 101.5000 150.9600 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8396 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.037 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.4668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 46.8448 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 242.82 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 102.2800 150.4750 102.4200 150.9600 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0518 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.4278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 66.752 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 54.2279 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 289.915 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 102.7400 150.4750 102.8800 150.9600 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6343 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.9455 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 29.4869 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 144.925 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 103.6600 150.4750 103.8000 150.9600 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5839 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.6935 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 27.9087 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 137.034 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 104.5800 150.4750 104.7200 150.9600 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 5.72444 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.204 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 105.0400 150.4750 105.1800 150.9600 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7929 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.7385 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 25.4424 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 124.703 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 105.9600 150.4750 106.1000 150.9600 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7307 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.3095 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 28.3046 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 137.628 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 106.8800 150.4750 107.0200 150.9600 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5586 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.632 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.8668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.76 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 50.8388 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 261.709 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 107.3400 150.4750 107.4800 150.9600 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.731 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.127 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.3278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.552 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 25.5459 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 136.618 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 108.2600 150.4750 108.4000 150.9600 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.486 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.6848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 73.456 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 59.4238 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 318.354 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 109.1800 150.4750 109.3200 150.9600 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6931 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.2395 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 29.4077 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 140.485 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 109.6400 150.4750 109.7800 150.9600 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.986 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.9148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 26.619 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 140.675 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 110.5600 150.4750 110.7000 150.9600 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2011 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.7795 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 17.8194 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 86.8606 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 111.4800 150.4750 111.6200 150.9600 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8195 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.8715 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 25.1002 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 120.428 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 111.9400 150.4750 112.0800 150.9600 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0267 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.9075 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 27.4279 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 134.63 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 112.8600 150.4750 113.0000 150.9600 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5405 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.4765 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 30.4061 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 149.521 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 113.7800 150.4750 113.9200 150.9600 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.0755 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 27.0554 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 129.931 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 114.2400 150.4750 114.3800 150.9600 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.498 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.329 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.2628 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.872 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 73.7737 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 380.954 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 115.1600 150.4750 115.3000 150.9600 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.984 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.0288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.624 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 70.6852 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 366.404 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 116.0800 150.4750 116.2200 150.9600 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7071 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.3095 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 30.177 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 148.376 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 116.5400 150.4750 116.6800 150.9600 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8671 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.1095 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 25.5329 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 125.156 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 117.4600 150.4750 117.6000 150.9600 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.9045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 31.4384 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 154.683 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 118.3800 150.4750 118.5200 150.9600 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0899 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2235 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 11.6461 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 55.7212 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 118.8400 150.4750 118.9800 150.9600 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8401 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.9745 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 33.2994 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 163.988 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 119.7600 150.4750 119.9000 150.9600 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0267 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.9075 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 25.3972 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 124.477 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 120.6800 150.4750 120.8200 150.9600 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2019 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7835 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.74182 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.4727 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 121.6000 150.4750 121.7400 150.9600 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3935 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.7415 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 27.1859 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 131.749 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 122.0600 150.4750 122.2000 150.9600 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5671 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.6095 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 27.379 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 134.659 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 122.9800 150.4750 123.1200 150.9600 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3135 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.3415 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 14.2331 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 68.9293 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 123.9000 150.4750 124.0400 150.9600 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.9675 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 34.1034 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 165.172 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 124.3600 150.4750 124.5000 150.9600 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.695 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.314 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.7068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 52.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 42.2638 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 226.242 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 125.2800 150.4750 125.4200 150.9600 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.2000 150.4750 126.3400 150.9600 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.6600 150.4750 126.8000 150.9600 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.5800 150.4750 127.7200 150.9600 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.5000 150.4750 128.6400 150.9600 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.9600 150.4750 129.1000 150.9600 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.8800 150.4750 130.0200 150.9600 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.8000 150.4750 130.9400 150.9600 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.2600 150.4750 131.4000 150.9600 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.1800 150.4750 132.3200 150.9600 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.1000 150.4750 133.2400 150.9600 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.5600 150.4750 133.7000 150.9600 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.4800 150.4750 134.6200 150.9600 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.4000 150.4750 135.5400 150.9600 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.8600 150.4750 136.0000 150.9600 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.7800 150.4750 136.9200 150.9600 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.7000 150.4750 137.8400 150.9600 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.1600 150.4750 138.3000 150.9600 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.0800 150.4750 139.2200 150.9600 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.0000 150.4750 140.1400 150.9600 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.4600 150.4750 140.6000 150.9600 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.3800 150.4750 141.5200 150.9600 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.3000 150.4750 142.4400 150.9600 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.7600 150.4750 142.9000 150.9600 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.6800 150.4750 143.8200 150.9600 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.6000 150.4750 144.7400 150.9600 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.0600 150.4750 145.2000 150.9600 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.9800 150.4750 146.1200 150.9600 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.9000 150.4750 147.0400 150.9600 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.3600 150.4750 147.5000 150.9600 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.2800 150.4750 148.4200 150.9600 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.2000 150.4750 149.3400 150.9600 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.1200 150.4750 150.2600 150.9600 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.1200 0.0000 150.2600 0.4850 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.2000 0.0000 149.3400 0.4850 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.8200 0.0000 147.9600 0.4850 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.4400 0.0000 146.5800 0.4850 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.0600 0.0000 145.2000 0.4850 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.6800 0.0000 143.8200 0.4850 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.3000 0.0000 142.4400 0.4850 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.9200 0.0000 141.0600 0.4850 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.5400 0.0000 139.6800 0.4850 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.6200 0.0000 138.7600 0.4850 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.2400 0.0000 137.3800 0.4850 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.8600 0.0000 136.0000 0.4850 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.4800 0.0000 134.6200 0.4850 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.1000 0.0000 133.2400 0.4850 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.7200 0.0000 131.8600 0.4850 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.3400 0.0000 130.4800 0.4850 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.9600 0.0000 129.1000 0.4850 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.0400 0.0000 128.1800 0.4850 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.6600 0.0000 126.8000 0.4850 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.2800 0.0000 125.4200 0.4850 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.9000 0.0000 124.0400 0.4850 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.5200 0.0000 122.6600 0.4850 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.1400 0.0000 121.2800 0.4850 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.7600 0.0000 119.9000 0.4850 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.3800 0.0000 118.5200 0.4850 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.4600 0.0000 117.6000 0.4850 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.0800 0.0000 116.2200 0.4850 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.7000 0.0000 114.8400 0.4850 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.3200 0.0000 113.4600 0.4850 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.9400 0.0000 112.0800 0.4850 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.5600 0.0000 110.7000 0.4850 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.1800 0.0000 109.3200 0.4850 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.8000 0.0000 107.9400 0.4850 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.8800 0.0000 107.0200 0.4850 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.5000 0.0000 105.6400 0.4850 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.1200 0.0000 104.2600 0.4850 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.7400 0.0000 102.8800 0.4850 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.3600 0.0000 101.5000 0.4850 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.8743 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.2635 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.9800 0.0000 100.1200 0.4850 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.7455 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.6195 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 98.6000 0.0000 98.7400 0.4850 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.9021 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.2845 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 97.2200 0.0000 97.3600 0.4850 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.2551 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.1675 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 96.3000 0.0000 96.4400 0.4850 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2255 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 94.9200 0.0000 95.0600 0.4850 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.7497 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.6405 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 93.5400 0.0000 93.6800 0.4850 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.578 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.536 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 10.5926 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 52.3929 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 92.1600 0.0000 92.3000 0.4850 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0508 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.74 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 36.3376 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 176.063 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.498027 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 36.9027 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 180.135 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.588117 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 40.7351 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 202.694 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.588117 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 90.7800 0.0000 90.9200 0.4850 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.43 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.989 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.217 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.2948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 29.9432 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 160.757 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 89.4000 0.0000 89.5400 0.4850 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4776 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.109 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.3778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 61.152 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 25.6257 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 137.73 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 88.0200 0.0000 88.1600 0.4850 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5345 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3185 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 3.45608 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 16.4831 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 86.6400 0.0000 86.7800 0.4850 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.2156 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.607 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.9474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.296 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met3  ;
    ANTENNAMAXAREACAR 18.3676 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 95.3365 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.538994 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.2916 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.496 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 52.8082 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 281.138 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.538994 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 85.7200 0.0000 85.8600 0.4850 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9176 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.427 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.672 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 4.30811 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 24.036 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 84.3400 0.0000 84.4800 0.4850 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6008 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.843 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.894 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.2936 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 119.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 50.2108 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 269.91 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 82.9600 0.0000 83.1000 0.4850 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0388 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.033 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.214 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.0316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 171.296 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 72.1432 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 385.802 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 81.5800 0.0000 81.7200 0.4850 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6224 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.725 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 59.6929 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 286.175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 62.3198 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 303.889 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.1468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 59.92 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 87.4252 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 438.844 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 80.2000 0.0000 80.3400 0.4850 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1494 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.468 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.7166 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.096 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 30.8932 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 166.883 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 78.8200 0.0000 78.9600 0.4850 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2172 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.1786 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.36 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 38.8454 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 196.588 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.678207 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.5238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.264 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 60.2954 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 312.048 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.678207 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 77.4400 0.0000 77.5800 0.4850 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 22.2426 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 110.6 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 194.207 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 956.952 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.0426 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.352 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 305.656 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1554.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.8646 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 85.552 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 341.387 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1747.67 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 76.0600 0.0000 76.2000 0.4850 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5192 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.1069 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.032 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 168.088 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 871.702 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.8057 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 106.096 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 212.696 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1110.66 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 75.1400 0.0000 75.2800 0.4850 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.967 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.5319 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.9854 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 140 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 58.5257 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 315.315 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 73.7600 0.0000 73.9000 0.4850 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.685 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 77.9079 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 386.389 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.31746 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 79.9317 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 400.738 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.634921 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.6348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.856 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 101.632 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 517.531 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.634921 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 72.3800 0.0000 72.5200 0.4850 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.873 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.1749 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 154.555 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 798.925 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.8706 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 197.584 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 237.597 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1243.93 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 71.0000 0.0000 71.1400 0.4850 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.43 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.989 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.527 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.9366 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 85.936 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 35.8932 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 193.55 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 69.6200 0.0000 69.7600 0.4850 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.4297 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.6865 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 21.2381 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 105.15 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 68.2400 0.0000 68.3800 0.4850 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.6009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 77.5425 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 35.1372 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 174.645 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 66.8600 0.0000 67.0000 0.4850 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1986 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.832 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.7657 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 182.312 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 956.75 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.9097 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 191.984 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 263.19 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1389.15 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 65.4800 0.0000 65.6200 0.4850 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.2534 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.985 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 112.397 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 549.619 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.6507 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.936 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 134.133 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 666.592 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 64.5600 0.0000 64.7000 0.4850 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.1411 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 110.093 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 49.8673 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 247.956 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.0900901 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.7408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.088 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 56.0403 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 281.938 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0900901 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 63.1800 0.0000 63.3200 0.4850 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.4637 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.8665 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 23.5669 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 116.816 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 61.8000 0.0000 61.9400 0.4850 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0994 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.4945 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 206.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 86.6993 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 464.505 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 60.4200 0.0000 60.5600 0.4850 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.6625 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 87.9585 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 39.7804 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 198.105 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 59.0400 0.0000 59.1800 0.4850 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.056 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.6824 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 154.384 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 64.6 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 347.712 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 57.6600 0.0000 57.8000 0.4850 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.05 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.863 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 78.1484 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 378.452 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 80.2829 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 392.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.6568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 30.64 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 93.0235 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 462.001 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 56.2800 0.0000 56.4200 0.4850 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.5099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 91.9695 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 41.689 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 207.139 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 54.9000 0.0000 55.0400 0.4850 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.0036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.395 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 31.6137 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 147.565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.498027 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 32.3592 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 152.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.588117 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.2968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 108.72 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 78.0727 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 397.457 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.588117 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 53.9800 0.0000 54.1200 0.4850 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.9625 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.4685 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 26.9426 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 133.938 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 52.6000 0.0000 52.7400 0.4850 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5264 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.471 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.4633 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 206.544 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.109 LAYER met4  ;
    ANTENNAMAXAREACAR 34.6829 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 186.243 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 51.2200 0.0000 51.3600 0.4850 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.6383 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.0835 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 49.8400 0.0000 49.9800 0.4850 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.8693 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.0295 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.465 LAYER met2  ;
    ANTENNAMAXAREACAR 4.00268 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.6333 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.023088 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.3985 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.728 LAYER met3  ;
    ANTENNAGATEAREA 9.1575 LAYER met3  ;
    ANTENNAMAXAREACAR 4.5922 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 22.8796 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.023088 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 48.4600 0.0000 48.6000 0.4850 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.8791 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.1275 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.465 LAYER met2  ;
    ANTENNAMAXAREACAR 9.63016 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.0596 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.291371 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.3985 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.728 LAYER met3  ;
    ANTENNAGATEAREA 9.1575 LAYER met3  ;
    ANTENNAMAXAREACAR 10.7444 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 51.5453 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 47.0800 0.0000 47.2200 0.4850 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.8595 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.8825 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.465 LAYER met2  ;
    ANTENNAMAXAREACAR 3.99986 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.5909 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.023088 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.3985 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.728 LAYER met3  ;
    ANTENNAGATEAREA 9.1575 LAYER met3  ;
    ANTENNAMAXAREACAR 4.58937 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 22.8372 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.023088 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 45.7000 0.0000 45.8400 0.4850 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8487 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2335 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 44.3200 0.0000 44.4600 0.4850 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.3315 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 43.4000 0.0000 43.5400 0.4850 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 42.0200 0.0000 42.1600 0.4850 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 40.6400 0.0000 40.7800 0.4850 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 39.2600 0.0000 39.4000 0.4850 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 37.8800 0.0000 38.0200 0.4850 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 36.5000 0.0000 36.6400 0.4850 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 35.1200 0.0000 35.2600 0.4850 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.3315 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 33.7400 0.0000 33.8800 0.4850 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.3315 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 32.8200 0.0000 32.9600 0.4850 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 31.4400 0.0000 31.5800 0.4850 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 30.0600 0.0000 30.2000 0.4850 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 28.6800 0.0000 28.8200 0.4850 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 27.3000 0.0000 27.4400 0.4850 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 25.9200 0.0000 26.0600 0.4850 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 24.5400 0.0000 24.6800 0.4850 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.3315 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 23.1600 0.0000 23.3000 0.4850 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.3315 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 22.2400 0.0000 22.3800 0.4850 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 20.8600 0.0000 21.0000 0.4850 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 19.4800 0.0000 19.6200 0.4850 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 18.1000 0.0000 18.2400 0.4850 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 16.7200 0.0000 16.8600 0.4850 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 15.3400 0.0000 15.4800 0.4850 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 13.9600 0.0000 14.1000 0.4850 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.3315 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 12.5800 0.0000 12.7200 0.4850 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.3315 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 11.6600 0.0000 11.8000 0.4850 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 10.2800 0.0000 10.4200 0.4850 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 8.9000 0.0000 9.0400 0.4850 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 7.5200 0.0000 7.6600 0.4850 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 6.1400 0.0000 6.2800 0.4850 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 4.7600 0.0000 4.9000 0.4850 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.2825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 3.3800 0.0000 3.5200 0.4850 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.3315 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2.0000 0.0000 2.1400 0.4850 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8389 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.0865 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1.0800 0.0000 1.2200 0.4850 ;
    END
  END io_oeb[0]
  PIN irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1413 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5985 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 148.3400 0.4850 148.4800 ;
    END
  END irq[2]
  PIN irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 149.0200 0.4850 149.1600 ;
    END
  END irq[1]
  PIN irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.5256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.402 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 150.0400 0.4850 150.1800 ;
    END
  END irq[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT 24.0200 24.1200 32.0200 126.8400 ;
        RECT 118.8600 24.1200 126.8600 126.8400 ;
        RECT 40.8000 24.1200 44.1600 126.8400 ;
        RECT 68.0000 24.1200 71.3600 126.8400 ;
        RECT 95.2000 24.1200 98.5600 126.8400 ;
      LAYER met5 ;
        RECT 24.0200 24.1200 126.8600 32.1200 ;
        RECT 24.0200 40.8000 126.8600 44.1600 ;
        RECT 24.0200 68.0000 126.8600 71.3600 ;
        RECT 24.0200 118.8400 126.8600 126.8400 ;
        RECT 24.0200 95.2000 126.8600 98.5600 ;
    END
# end of P/G power stripe data as pin

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT 8.0200 8.1200 16.0200 142.8400 ;
        RECT 134.8600 8.1200 142.8600 142.8400 ;
        RECT 54.4000 8.1200 57.7600 142.8400 ;
        RECT 81.6000 8.1200 84.9600 142.8400 ;
        RECT 27.2000 8.1200 30.5600 11.4800 ;
      LAYER met5 ;
        RECT 8.0200 8.1200 142.8600 16.1200 ;
        RECT 8.0200 54.4000 142.8600 57.7600 ;
        RECT 8.0200 27.2000 11.3800 30.5600 ;
        RECT 8.0200 134.8400 142.8600 142.8400 ;
        RECT 8.0200 81.6000 142.8600 84.9600 ;
    END
# end of P/G power stripe data as pin

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.0000 0.0000 150.8800 150.9600 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 150.8800 150.9600 ;
    LAYER met2 ;
      RECT 0.0000 0.0000 150.8800 150.9600 ;
    LAYER met3 ;
      RECT 0.0000 0.0000 150.8800 150.9600 ;
    LAYER met4 ;
      RECT 0.0000 0.0000 150.8800 150.9600 ;
    LAYER met5 ;
      RECT 0.0000 0.0000 150.8800 150.9600 ;
  END
END user_proj_example

END LIBRARY
