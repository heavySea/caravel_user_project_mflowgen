##
## LEF for PtnCells ;
## created by Innovus v17.11-s080_1 on Thu Jun 17 18:21:47 2021
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO user_proj_example
  CLASS BLOCK ;
  SIZE 150.8800 BY 150.9600 ;
  FOREIGN user_proj_example 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 23.1126 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 124.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.492 LAYER met4  ;
    ANTENNAMAXAREACAR 49.5944 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 261.437 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.267073 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 150.0400 150.8800 150.1800 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.623 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 41.8623 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 203.135 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 148.6800 150.8800 148.8200 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5416 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.482 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 56.506 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 271.679 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 147.3200 150.8800 147.4600 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7789 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.6685 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 47.5048 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 233.214 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 145.9600 150.8800 146.1000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6025 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.7865 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.504 LAYER met2  ;
    ANTENNAMAXAREACAR 32.1514 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 150.689 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 144.6000 150.8800 144.7400 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3605 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 53.9321 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 262.262 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 143.2400 150.8800 143.3800 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8185 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.8665 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 40.6091 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 195.54 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 141.5400 150.8800 141.6800 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 50.9377 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 247.29 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 140.1800 150.8800 140.3200 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2527 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.5003 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 23.1258 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 124.683 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 138.8200 150.8800 138.9600 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3235 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 6.22485 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.2606 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 137.4600 150.8800 137.6000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.623 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 26.0903 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 127.915 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 136.1000 150.8800 136.2400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.8755 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.0985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.1648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 35.0438 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 184.947 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 134.7400 150.8800 134.8800 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 25.519 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 125.059 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 133.0400 150.8800 133.1800 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 25.2588 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 123.758 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 131.6800 150.8800 131.8200 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.623 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 24.6648 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 120.788 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 130.3200 150.8800 130.4600 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4188 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.868 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 18.8152 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 91.303 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 128.9600 150.8800 129.1000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.887 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.973 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 24.902 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 120.166 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 127.6000 150.8800 127.7400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.2045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.4438 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 38.696 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 204.111 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 125.9000 150.8800 126.0400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7956 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.752 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 5.31697 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.7212 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 124.5400 150.8800 124.6800 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3493 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.9488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.864 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 12.0131 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 64.103 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 123.1800 150.8800 123.3200 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0714 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.225 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 119 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.8658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.088 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 46.4333 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 248.251 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 121.8200 150.8800 121.9600 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1995 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.394 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.8834 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 59.456 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 51.3941 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 277.299 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 120.4600 150.8800 120.6000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.437 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.0458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.256 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 58.864 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 92.136 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met5  ;
    ANTENNAMAXAREACAR 250.671 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 424.038 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 119.1000 150.8800 119.2400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4439 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 14.0588 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 73.1818 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 117.4000 150.8800 117.5400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.217 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.924 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.2158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.496 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 93.088 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 143.472 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 147.093 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 243.203 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 116.0400 150.8800 116.1800 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3303 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.4258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.408 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 34.1246 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 181.56 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 114.6800 150.8800 114.8200 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.161 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 148.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.8846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.992 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 12.2911 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 68.0404 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 113.3200 150.8800 113.4600 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.469 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.8718 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.92 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 5.04667 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 27.9636 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 111.9600 150.8800 112.1000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.161 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.871 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.2878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.88 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 52.24 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 82.2 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met5  ;
    ANTENNAMAXAREACAR 236.004 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 447.101 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 110.2600 150.8800 110.4000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1022 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.45345 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 135.712 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 207.408 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 213.205 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 355.605 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 108.9000 150.8800 109.0400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.4835 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.1385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.97 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 117.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.6698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 37.081 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 196.98 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 107.5400 150.8800 107.6800 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1645 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.4838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.592 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 41.2 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 65.64 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met5  ;
    ANTENNAMAXAREACAR 197.106 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 411.747 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 106.1800 150.8800 106.3200 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1449 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.1678 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 145.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 7.48303 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 39.7657 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 104.8200 150.8800 104.9600 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.609 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.8758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 49.016 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 91.888 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 141.672 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 145.564 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 241.26 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 103.4600 150.8800 103.6000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.3248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.744 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 136.144 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 208.056 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 209.147 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 332.089 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 101.7600 150.8800 101.9000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4213 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.8275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.0608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.128 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 30.7453 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 162.586 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 100.4000 150.8800 100.5400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9755 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.225 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 119 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.1818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 49.44 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 44.5642 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 237.055 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 99.0400 150.8800 99.1800 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5576 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.562 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 3.21434 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.299 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 97.6800 150.8800 97.8200 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.4708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.856 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 142 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 216.84 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 218.267 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 346.57 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 96.3200 150.8800 96.4600 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.4365 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 32.0406 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 156.863 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 94.6200 150.8800 94.7600 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3691 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6195 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 19.8176 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 96.2242 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 93.2600 150.8800 93.4000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 91.9000 150.8800 92.0400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 90.5400 150.8800 90.6800 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 89.1800 150.8800 89.3200 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 87.8200 150.8800 87.9600 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 86.1200 150.8800 86.2600 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 84.7600 150.8800 84.9000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 83.4000 150.8800 83.5400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 82.0400 150.8800 82.1800 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 80.6800 150.8800 80.8200 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 78.9800 150.8800 79.1200 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 77.6200 150.8800 77.7600 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 76.2600 150.8800 76.4000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 74.9000 150.8800 75.0400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 73.5400 150.8800 73.6800 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 72.1800 150.8800 72.3200 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 70.4800 150.8800 70.6200 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 69.1200 150.8800 69.2600 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 67.7600 150.8800 67.9000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 66.4000 150.8800 66.5400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 65.0400 150.8800 65.1800 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 63.3400 150.8800 63.4800 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 61.9800 150.8800 62.1200 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 60.6200 150.8800 60.7600 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 59.2600 150.8800 59.4000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 57.9000 150.8800 58.0400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 56.5400 150.8800 56.6800 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 54.8400 150.8800 54.9800 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 53.4800 150.8800 53.6200 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 52.1200 150.8800 52.2600 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 50.7600 150.8800 50.9000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 49.4000 150.8800 49.5400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3950 47.7000 150.8800 47.8400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4144 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.846 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 30.5623 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 142.409 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 46.3400 150.8800 46.4800 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0658 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.9728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.992 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 44.9800 150.8800 45.1200 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8623 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.0325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.2358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.728 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 43.6200 150.8800 43.7600 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 42.2600 150.8800 42.4000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.2132 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.84 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 40.9000 150.8800 41.0400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.8203 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.9935 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 39.2000 150.8800 39.3400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.1733 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.6405 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 37.8400 150.8800 37.9800 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 36.4800 150.8800 36.6200 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.5437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.4395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.7468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.12 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 35.1200 150.8800 35.2600 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.046 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.886 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 33.7600 150.8800 33.9000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0966 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.292 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 98.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.9638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.944 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 32.0600 150.8800 32.2000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 30.7000 150.8800 30.8400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 29.3400 150.8800 29.4800 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 27.9800 150.8800 28.1200 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 26.6200 150.8800 26.7600 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.842 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.984 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 25.2600 150.8800 25.4000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7665 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.5535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.5048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.496 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 23.5600 150.8800 23.7000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.969 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.619 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 22.2000 150.8800 22.3400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.2648 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.098 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 20.8400 150.8800 20.9800 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0156 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.852 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 19.4800 150.8800 19.6200 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.0908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.228 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 18.1200 150.8800 18.2600 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1372 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.46 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 16.4200 150.8800 16.5600 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.738 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.529 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.8388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.944 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 15.0600 150.8800 15.2000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 13.7000 150.8800 13.8400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.2505 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 12.3400 150.8800 12.4800 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.1429 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.4885 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 10.9800 150.8800 11.1200 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.2476 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.012 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 9.6200 150.8800 9.7600 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.39 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.724 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 7.9200 150.8800 8.0600 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.8489 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.0185 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 6.5600 150.8800 6.7000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.2465 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.0065 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 5.2000 150.8800 5.3400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.04 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.974 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 3.8400 150.8800 3.9800 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.6417 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.9825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 2.4800 150.8800 2.6200 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1204 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.376 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 150.3950 1.1200 150.8800 1.2600 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 0.7800 0.4850 0.9200 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 1.4600 0.4850 1.6000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 2.1400 0.4850 2.2800 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 2.8200 0.4850 2.9600 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 3.8400 0.4850 3.9800 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 4.5200 0.4850 4.6600 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 5.2000 0.4850 5.3400 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 6.2200 0.4850 6.3600 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 6.9000 0.4850 7.0400 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 7.5800 0.4850 7.7200 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 8.2600 0.4850 8.4000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 9.2800 0.4850 9.4200 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 9.9600 0.4850 10.1000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 10.6400 0.4850 10.7800 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 11.6600 0.4850 11.8000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 12.3400 0.4850 12.4800 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 13.0200 0.4850 13.1600 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 14.0400 0.4850 14.1800 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 14.7200 0.4850 14.8600 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 15.4000 0.4850 15.5400 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 16.0800 0.4850 16.2200 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 17.1000 0.4850 17.2400 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 17.7800 0.4850 17.9200 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 18.4600 0.4850 18.6000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 19.4800 0.4850 19.6200 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.1600 0.4850 20.3000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.8400 0.4850 20.9800 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 21.8600 0.4850 22.0000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 22.5400 0.4850 22.6800 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 23.2200 0.4850 23.3600 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 23.9000 0.4850 24.0400 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 24.9200 0.4850 25.0600 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 25.6000 0.4850 25.7400 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 26.2800 0.4850 26.4200 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 27.3000 0.4850 27.4400 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 27.9800 0.4850 28.1200 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 28.6600 0.4850 28.8000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 29.6800 0.4850 29.8200 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 30.3600 0.4850 30.5000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 31.0400 0.4850 31.1800 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 31.7200 0.4850 31.8600 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 32.7400 0.4850 32.8800 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 33.4200 0.4850 33.5600 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 34.1000 0.4850 34.2400 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 35.1200 0.4850 35.2600 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 35.8000 0.4850 35.9400 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 36.4800 0.4850 36.6200 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 37.5000 0.4850 37.6400 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 38.1800 0.4850 38.3200 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 38.8600 0.4850 39.0000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 39.5400 0.4850 39.6800 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 40.5600 0.4850 40.7000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 41.2400 0.4850 41.3800 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 41.9200 0.4850 42.0600 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 42.9400 0.4850 43.0800 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 43.6200 0.4850 43.7600 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 44.3000 0.4850 44.4400 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 45.3200 0.4850 45.4600 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 46.0000 0.4850 46.1400 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 46.6800 0.4850 46.8200 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 47.3600 0.4850 47.5000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 48.3800 0.4850 48.5200 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2225 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 7.66824 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 26.0189 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 49.0600 0.4850 49.2000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6848 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.263 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.6828 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 132.112 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.492 LAYER met3  ;
    ANTENNAMAXAREACAR 52.0468 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 276.702 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.185772 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 49.7400 0.4850 49.8800 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6858 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.085 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 36.303 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 177.881 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 50.7600 0.4850 50.9000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0994 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.8088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.784 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 49.6036 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 247.596 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 51.4400 0.4850 51.5800 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2096 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.822 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 74.5212 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 369.299 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 52.1200 0.4850 52.2600 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 94.7396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 358.03 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 52.8000 0.4850 52.9400 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0641 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.632 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 158.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.3798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 65.2976 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 348.408 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 53.8200 0.4850 53.9600 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8052 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.8 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 23.6784 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 115.234 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 54.5000 0.4850 54.6400 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.301 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.344 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.307 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 146.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 17.4436 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 91.6687 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 55.1800 0.4850 55.3200 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2353 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.605 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 126.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.4868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.4 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 36.0699 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 190.174 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 56.2000 0.4850 56.3400 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0854 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.755 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 143.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.1656 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.824 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 15.8335 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 86.6424 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 56.8800 0.4850 57.0200 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1232 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.45345 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 132.064 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 201.936 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 214.448 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 388.347 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 57.5600 0.4850 57.7000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2478 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.078 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.7778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.16 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 76.528 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 118.632 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 141.855 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 315.21 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 58.5800 0.4850 58.7200 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.854 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.2428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.432 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 38.3053 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 199.673 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 59.2600 0.4850 59.4000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6781 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.8426 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.44 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 71.008 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 110.352 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 119.824 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 221.575 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 59.9400 0.4850 60.0800 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3892 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.806 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3924 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.776 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 41.2 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 65.64 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met5  ;
    ANTENNAMAXAREACAR 202.8 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 440.836 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 60.6200 0.4850 60.7600 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 46.4501 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 229.271 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 61.6400 0.4850 61.7800 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9755 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.1098 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 63.5446 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 335.919 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 62.3200 0.4850 62.4600 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.091 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.2838 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.984 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 85.88 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 452.513 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 63.0000 0.4850 63.1400 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.0168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.56 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 18.836 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 97.196 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 64.0200 0.4850 64.1600 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.672 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.199 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.338 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 8.60444 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 48.501 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 64.7000 0.4850 64.8400 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0742 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.2474 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 39.7584 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 216.057 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 65.3800 0.4850 65.5200 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6525 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.0988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.664 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 59.8533 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 317.22 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 66.4000 0.4850 66.5400 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.83 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.3668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.76 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 77.5931 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 404.933 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 67.0800 0.4850 67.2200 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.161 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.525 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.7998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.944 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 98.608 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 151.752 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 152.682 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 240.832 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 67.7600 0.4850 67.9000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1372 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.4226 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.528 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 70.0392 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 371.624 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 68.4400 0.4850 68.5800 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2152 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.896 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 14.6493 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 74.4162 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 69.4600 0.4850 69.6000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 27.1976 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 133.307 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 70.1400 0.4850 70.2800 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9255 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.4328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.112 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 40.8788 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 213.37 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 70.8200 0.4850 70.9600 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 24.556 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 120.099 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 71.8400 0.4850 71.9800 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1413 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5985 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 27.4192 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 130.428 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 72.5200 0.4850 72.6600 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 32.9616 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 162.127 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 73.2000 0.4850 73.3400 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5121 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3345 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 7.44121 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.0485 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 74.2200 0.4850 74.3600 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9492 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.3288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 98.224 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 76.8012 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 406.501 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 74.9000 0.4850 75.0400 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 75.5800 0.4850 75.7200 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 76.2600 0.4850 76.4000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 77.2800 0.4850 77.4200 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 77.9600 0.4850 78.1000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 78.6400 0.4850 78.7800 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 79.6600 0.4850 79.8000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 80.3400 0.4850 80.4800 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 81.0200 0.4850 81.1600 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 82.0400 0.4850 82.1800 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 82.7200 0.4850 82.8600 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 83.4000 0.4850 83.5400 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 84.0800 0.4850 84.2200 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 85.1000 0.4850 85.2400 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 85.7800 0.4850 85.9200 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 86.4600 0.4850 86.6000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 87.4800 0.4850 87.6200 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 88.1600 0.4850 88.3000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 88.8400 0.4850 88.9800 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 89.8600 0.4850 90.0000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 90.5400 0.4850 90.6800 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 91.2200 0.4850 91.3600 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 91.9000 0.4850 92.0400 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 92.9200 0.4850 93.0600 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 93.6000 0.4850 93.7400 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 94.2800 0.4850 94.4200 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 95.3000 0.4850 95.4400 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 95.9800 0.4850 96.1200 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 96.6600 0.4850 96.8000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 97.6800 0.4850 97.8200 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 98.3600 0.4850 98.5000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 99.0400 0.4850 99.1800 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.0000 99.7200 0.4850 99.8600 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 100.7400 0.4850 100.8800 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0882 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.8618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.4 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 101.4200 0.4850 101.5600 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 102.1000 0.4850 102.2400 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3605 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 103.1200 0.4850 103.2600 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 103.8000 0.4850 103.9400 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.176 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.654 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 104.4800 0.4850 104.6200 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 105.1600 0.4850 105.3000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4417 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 106.1800 0.4850 106.3200 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 106.8600 0.4850 107.0000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.5028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.288 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 107.5400 0.4850 107.6800 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0497 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.3848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.856 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 108.5600 0.4850 108.7000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 109.2400 0.4850 109.3800 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 109.9200 0.4850 110.0600 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1889 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8365 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 110.9400 0.4850 111.0800 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 111.6200 0.4850 111.7600 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8954 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.133 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 112.3000 0.4850 112.4400 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0798 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.2968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.72 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 112.9800 0.4850 113.1200 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8432 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.99 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 114.0000 0.4850 114.1400 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3314 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.431 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 114.6800 0.4850 114.8200 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 115.3600 0.4850 115.5000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9268 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.473 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.3988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.264 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 116.3800 0.4850 116.5200 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 117.0600 0.4850 117.2000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.9951 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.8675 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 117.7400 0.4850 117.8800 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.542 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.484 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 118.7600 0.4850 118.9000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3304 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.491 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.0528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.752 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 119.4400 0.4850 119.5800 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3524 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.536 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 120.1200 0.4850 120.2600 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9422 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.485 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 120.8000 0.4850 120.9400 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1722 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.1358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.528 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 121.8200 0.4850 121.9600 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0332 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 122.5000 0.4850 122.6400 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8592 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.07 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 123.1800 0.4850 123.3200 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 124.2000 0.4850 124.3400 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1004 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.223 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.3658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.088 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 124.8800 0.4850 125.0200 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3031 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.2365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.9258 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.408 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 125.5600 0.4850 125.7000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 126.5800 0.4850 126.7200 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0854 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.898 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.1578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.312 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 127.2600 0.4850 127.4000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 127.9400 0.4850 128.0800 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8984 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.266 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 128.6200 0.4850 128.7600 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 129.6400 0.4850 129.7800 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.0548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.096 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 130.3200 0.4850 130.4600 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3672 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.61 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 131.0000 0.4850 131.1400 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5721 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.5815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.3298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.896 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 132.0200 0.4850 132.1600 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 132.7000 0.4850 132.8400 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3588 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.568 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 133.3800 0.4850 133.5200 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.5956 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.752 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 134.4000 0.4850 134.5400 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.898 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.264 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 135.0800 0.4850 135.2200 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0966 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.887 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.7328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 57.712 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 135.7600 0.4850 135.9000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2779 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.752 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.3298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 60.896 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 136.4400 0.4850 136.5800 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1498 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.47 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.2508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.808 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 137.4600 0.4850 137.6000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6052 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 138.1400 0.4850 138.2800 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0324 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.936 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 138.8200 0.4850 138.9600 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.6897 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.2225 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 139.8400 0.4850 139.9800 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.3605 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 140.5200 0.4850 140.6600 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3668 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.673 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.5018 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.48 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 141.2000 0.4850 141.3400 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.2864 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.206 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 142.2200 0.4850 142.3600 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6129 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8385 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 142.9000 0.4850 143.0400 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.2711 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.2475 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 143.5800 0.4850 143.7200 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1413 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5985 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 144.2600 0.4850 144.4000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0714 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.1785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.287 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.3668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 55.76 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 145.2800 0.4850 145.4200 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8763 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.1555 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 145.9600 0.4850 146.1000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3199 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.2228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.992 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 146.6400 0.4850 146.7800 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1504 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.644 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 147.6600 0.4850 147.8000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0685 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2345 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.6200 150.4750 0.7600 150.9600 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8427 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1055 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1.0800 150.4750 1.2200 150.9600 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1316 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.497 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.189 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.0748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.536 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2.0000 150.4750 2.1400 150.9600 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.62 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.9288 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 69.424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2.9200 150.4750 3.0600 150.9600 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.351 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.9788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 91.024 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 3.3800 150.4750 3.5200 150.9600 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.3763 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.6555 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 4.3000 150.4750 4.4400 150.9600 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.3963 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.7555 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 5.2200 150.4750 5.3600 150.9600 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.6631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.0895 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 5.6800 150.4750 5.8200 150.9600 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4395 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 6.6000 150.4750 6.7400 150.9600 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2499 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0235 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 7.5200 150.4750 7.6600 150.9600 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.6902 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.29 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.2288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.024 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 7.9800 150.4750 8.1200 150.9600 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.8671 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.1095 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 8.9000 150.4750 9.0400 150.9600 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.2647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.0975 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 9.8200 150.4750 9.9600 150.9600 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.8219 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.8835 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 10.2800 150.4750 10.4200 150.9600 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0643 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2135 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 11.2000 150.4750 11.3400 150.9600 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.5027 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.2875 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 12.1200 150.4750 12.2600 150.9600 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.698 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.7328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.712 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 12.5800 150.4750 12.7200 150.9600 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6224 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.833 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.1088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.384 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 13.5000 150.4750 13.6400 150.9600 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.2842 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.26 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.4428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.832 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 14.4200 150.4750 14.5600 150.9600 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0384 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 14.8800 150.4750 15.0200 150.9600 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3283 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4155 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 15.8000 150.4750 15.9400 150.9600 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.8575 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.1795 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 16.7200 150.4750 16.8600 150.9600 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.1821 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.5665 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 17.1800 150.4750 17.3200 150.9600 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.6495 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.1395 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 18.1000 150.4750 18.2400 150.9600 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.664 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.1928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.832 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 19.0200 150.4750 19.1600 150.9600 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6355 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0695 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 19.4800 150.4750 19.6200 150.9600 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.2003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.7755 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 20.4000 150.4750 20.5400 150.9600 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.487 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.274 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.712 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.3538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 45.024 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 21.3200 150.4750 21.4600 150.9600 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4635 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 21.7800 150.4750 21.9200 150.9600 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7723 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.6355 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 22.7000 150.4750 22.8400 150.9600 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.5503 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.5255 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 23.6200 150.4750 23.7600 150.9600 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.2811 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.1795 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 24.0800 150.4750 24.2200 150.9600 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0643 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2135 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 25.0000 150.4750 25.1400 150.9600 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.2215 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.9995 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 25.9200 150.4750 26.0600 150.9600 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.6599 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.0735 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 26.3800 150.4750 26.5200 150.9600 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.591 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.794 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.513 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.6376 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 159.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 66.4978 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 342.159 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.844157 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 27.3000 150.4750 27.4400 150.9600 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.772 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.578 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.031 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.5786 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 185.36 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 118.261 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 614.673 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.946868 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 28.2200 150.4750 28.3600 150.9600 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.514 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 71.5479 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 352.208 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 28.6800 150.4750 28.8200 150.9600 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4776 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.7698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 84.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 35.5176 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 190.486 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 29.6000 150.4750 29.7400 150.9600 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.6848 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.06 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 27.453 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 126.762 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 30.5200 150.4750 30.6600 150.9600 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1368 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.287 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 46.3893 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 226.687 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.287421 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.7468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.12 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 79.6028 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 404.885 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.287421 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 31.4400 150.4750 31.5800 150.9600 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.076 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 30.1915 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 144.987 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.358176 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.3096 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.592 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 44.4023 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 222.897 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 31.9000 150.4750 32.0400 150.9600 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5586 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.632 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.609 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.7356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 180.864 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 137.732 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 727.839 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.905577 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 32.8200 150.4750 32.9600 150.9600 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.3834 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.319 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 24.9715 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 119.16 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.498027 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 25.717 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 124.187 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.588117 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.6967 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 94.848 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 65.5744 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 337.809 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.588117 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 33.7400 150.4750 33.8800 150.9600 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.1764 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 85.603 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.6455 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 153.712 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 87.4605 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 457.881 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 34.2000 150.4750 34.3400 150.9600 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4846 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.262 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.375 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 103.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.8305 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 144.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 116.256 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 605.615 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.85635 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 35.1200 150.4750 35.2600 150.9600 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.2 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.9776 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 123.488 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 80.1341 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 425.12 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.538994 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 36.0400 150.4750 36.1800 150.9600 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.351 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.4376 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 88.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 37.0216 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 199.568 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 36.5000 150.4750 36.6400 150.9600 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.783 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.0841 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.5573 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 121.712 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 88.5103 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 464.043 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 37.4200 150.4750 37.5600 150.9600 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5018 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.348 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.4852 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.52 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 194.327 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1043.81 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.31746 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.4998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.136 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 215.723 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1158.98 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.413208 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 38.3400 150.4750 38.4800 150.9600 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.8276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.721 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 119.679 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 585.008 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.0188 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.904 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 135.487 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 670.377 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 38.8000 150.4750 38.9400 150.9600 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.779 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.734 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.911 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.2562 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 211.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 139.57 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 741.169 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 39.7200 150.4750 39.8600 150.9600 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.1872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.539 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 118.542 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 580.341 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.4668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.96 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 133.107 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 659.08 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 40.6400 150.4750 40.7800 150.9600 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.34 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.505 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.597 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 229.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 426.729 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2223.45 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 7.25317 LAYER via4  ;
    ANTENNADIFFAREA 0.429 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 48.928 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 77.232 LAYER met5  ;
    ANTENNAGATEAREA 0.444 LAYER met5  ;
    ANTENNAMAXAREACAR 536.927 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 2397.39 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 41.1000 150.4750 41.2400 150.9600 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.9383 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 94.2515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.3565 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 111.583 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 560.686 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 42.0200 150.4750 42.1600 150.9600 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.5698 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 117.334 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 208.318 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 1028.29 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.9848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.056 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 226.302 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1125.26 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 42.9400 150.4750 43.0800 150.9600 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8038 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.858 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.575 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.6837 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 100.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 45.538 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 239.893 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.413208 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 43.4000 150.4750 43.5400 150.9600 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.902 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.092 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.8857 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 175.856 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 104.346 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 551.921 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.413208 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 44.3200 150.4750 44.4600 150.9600 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.5143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 82.0365 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 134.967 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 661.369 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.135 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.52 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 143.975 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 713.115 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 147.539 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 733.187 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 45.2400 150.4750 45.3800 150.9600 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.351 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.1162 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 109.44 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.429 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 12.496 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 22.584 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met5  ;
    ANTENNAMAXAREACAR 28.1441 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 50.8649 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 45.7000 150.4750 45.8400 150.9600 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1564 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.621 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.1497 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 145.264 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 80.0634 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 424.052 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.413208 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 46.6200 150.4750 46.7600 150.9600 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.486 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.2716 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 157.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 125.784 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 657.277 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.905577 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 47.5400 150.4750 47.6800 150.9600 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.1572 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.648 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 80.1685 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 389.496 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.765079 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 48.0000 150.4750 48.1400 150.9600 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.3948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.836 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 36.3947 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 172.286 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.381392 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 48.9200 150.4750 49.0600 150.9600 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.8664 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.053 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.0868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 11.4568 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 62.1622 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 49.8400 150.4750 49.9800 150.9600 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.8542 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.992 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.3378 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.272 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 7.51757 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 41.1532 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 50.3000 150.4750 50.4400 150.9600 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6592 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.837 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.4878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 84.28 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.429 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 23.536 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 39.144 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.109 LAYER met5  ;
    ANTENNAMAXAREACAR 28.048 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 59.7819 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 51.2200 150.4750 51.3600 150.9600 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.1400 150.4750 52.2800 150.9600 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.6000 150.4750 52.7400 150.9600 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.5200 150.4750 53.6600 150.9600 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.4400 150.4750 54.5800 150.9600 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.9000 150.4750 55.0400 150.9600 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.8200 150.4750 55.9600 150.9600 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.7400 150.4750 56.8800 150.9600 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.2000 150.4750 57.3400 150.9600 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.1200 150.4750 58.2600 150.9600 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.0400 150.4750 59.1800 150.9600 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.5000 150.4750 59.6400 150.9600 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.4200 150.4750 60.5600 150.9600 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.3400 150.4750 61.4800 150.9600 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.2600 150.4750 62.4000 150.9600 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.7200 150.4750 62.8600 150.9600 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.6400 150.4750 63.7800 150.9600 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.5600 150.4750 64.7000 150.9600 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.0200 150.4750 65.1600 150.9600 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.9400 150.4750 66.0800 150.9600 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.8600 150.4750 67.0000 150.9600 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.3200 150.4750 67.4600 150.9600 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.2400 150.4750 68.3800 150.9600 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.1600 150.4750 69.3000 150.9600 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.6200 150.4750 69.7600 150.9600 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.5400 150.4750 70.6800 150.9600 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.4600 150.4750 71.6000 150.9600 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.9200 150.4750 72.0600 150.9600 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.8400 150.4750 72.9800 150.9600 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.7600 150.4750 73.9000 150.9600 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.2200 150.4750 74.3600 150.9600 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.1400 150.4750 75.2800 150.9600 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.0600 150.4750 76.2000 150.9600 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.5200 150.4750 76.6600 150.9600 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.4400 150.4750 77.5800 150.9600 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.3600 150.4750 78.5000 150.9600 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.8200 150.4750 78.9600 150.9600 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.7400 150.4750 79.8800 150.9600 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.6600 150.4750 80.8000 150.9600 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.1200 150.4750 81.2600 150.9600 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.0400 150.4750 82.1800 150.9600 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.9600 150.4750 83.1000 150.9600 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.4200 150.4750 83.5600 150.9600 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.3400 150.4750 84.4800 150.9600 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.2600 150.4750 85.4000 150.9600 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.7200 150.4750 85.8600 150.9600 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.6400 150.4750 86.7800 150.9600 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.5600 150.4750 87.7000 150.9600 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.0200 150.4750 88.1600 150.9600 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.9400 150.4750 89.0800 150.9600 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.8600 150.4750 90.0000 150.9600 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.7800 150.4750 90.9200 150.9600 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.2400 150.4750 91.3800 150.9600 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.1600 150.4750 92.3000 150.9600 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.0800 150.4750 93.2200 150.9600 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.5400 150.4750 93.6800 150.9600 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.4600 150.4750 94.6000 150.9600 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.3800 150.4750 95.5200 150.9600 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.8400 150.4750 95.9800 150.9600 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.7600 150.4750 96.9000 150.9600 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.6800 150.4750 97.8200 150.9600 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.1400 150.4750 98.2800 150.9600 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.0600 150.4750 99.2000 150.9600 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9643 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5955 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 5.30692 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.6478 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.161635 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 99.9800 150.4750 100.1200 150.9600 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4035 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.9095 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.665 LAYER met2  ;
    ANTENNAMAXAREACAR 10.4426 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 49.9804 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0772932 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 100.4400 150.4750 100.5800 150.9600 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6175 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.8615 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 27.7842 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 136.412 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 101.3600 150.4750 101.5000 150.9600 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5586 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.632 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.9148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 49.3972 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 254.089 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 102.2800 150.4750 102.4200 150.9600 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0941 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2445 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.84566 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.7596 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 102.7400 150.4750 102.8800 150.9600 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8586 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.014 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.4018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 45.28 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 50.4513 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 269.608 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 103.6600 150.4750 103.8000 150.9600 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8207 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8775 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 14.3895 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 69.4384 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 104.5800 150.4750 104.7200 150.9600 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2479 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.0135 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 26.0893 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 128.21 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 105.0400 150.4750 105.1800 150.9600 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.0975 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 33.0053 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 162.517 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 105.9600 150.4750 106.1000 150.9600 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6875 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 11.2804 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 54.1657 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 106.8800 150.4750 107.0200 150.9600 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0587 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.0675 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 18.2691 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 86.8929 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 107.3400 150.4750 107.4800 150.9600 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1079 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.3135 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 25.5236 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 125.382 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 108.2600 150.4750 108.4000 150.9600 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8687 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1175 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.6602 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.8828 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 109.1800 150.4750 109.3200 150.9600 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.4016 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.729 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.8788 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.824 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 13.8489 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 72.7354 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 109.6400 150.4750 109.7800 150.9600 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8979 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.2635 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 24.6752 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 121.139 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 110.5600 150.4750 110.7000 150.9600 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0427 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9875 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 5.05818 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.0545 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 111.4800 150.4750 111.6200 150.9600 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3123 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.3355 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 27.4053 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 134.517 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 111.9400 150.4750 112.0800 150.9600 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0267 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.9075 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 25.1956 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 123.741 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 112.8600 150.4750 113.0000 150.9600 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8979 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.2635 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 24.6752 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 121.139 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 113.7800 150.4750 113.9200 150.9600 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6931 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.2395 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 28.8315 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 138.812 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 114.2400 150.4750 114.3800 150.9600 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8569 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.0585 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 28.7515 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 141.248 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 115.1600 150.4750 115.3000 150.9600 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1219 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.3835 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 27.3042 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 131.176 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 116.0800 150.4750 116.2200 150.9600 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0923 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.2355 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 14.3216 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 69.099 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 116.5400 150.4750 116.6800 150.9600 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8695 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.1215 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 28.6008 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 140.768 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 117.4600 150.4750 117.6000 150.9600 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0001 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.7745 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 26.2796 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 128.889 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 118.3800 150.4750 118.5200 150.9600 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3424 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.551 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.0408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.688 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 45.6073 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 239.826 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 118.8400 150.4750 118.9800 150.9600 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1555 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.5515 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 25.9176 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 127.079 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 119.7600 150.4750 119.9000 150.9600 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0518 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.1928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.832 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 66.8489 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 347.859 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 120.6800 150.4750 120.8200 150.9600 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1595 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6895 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 20.0145 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 97.8909 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 121.6000 150.4750 121.7400 150.9600 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0477 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.0125 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 26.9923 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 132.453 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 122.0600 150.4750 122.2000 150.9600 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0025 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.7865 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 30.8889 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 149.992 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 122.9800 150.4750 123.1200 150.9600 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5363 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.4555 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 28.7063 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 141.022 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 123.9000 150.4750 124.0400 150.9600 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 7.43192 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.6505 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 124.3600 150.4750 124.5000 150.9600 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.8325 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 26.9527 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 132.255 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 125.2800 150.4750 125.4200 150.9600 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.2000 150.4750 126.3400 150.9600 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.6600 150.4750 126.8000 150.9600 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.5800 150.4750 127.7200 150.9600 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.5000 150.4750 128.6400 150.9600 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.9600 150.4750 129.1000 150.9600 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.8800 150.4750 130.0200 150.9600 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.8000 150.4750 130.9400 150.9600 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.2600 150.4750 131.4000 150.9600 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.1800 150.4750 132.3200 150.9600 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.1000 150.4750 133.2400 150.9600 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.5600 150.4750 133.7000 150.9600 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.4800 150.4750 134.6200 150.9600 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.4000 150.4750 135.5400 150.9600 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.8600 150.4750 136.0000 150.9600 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.7800 150.4750 136.9200 150.9600 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.7000 150.4750 137.8400 150.9600 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.1600 150.4750 138.3000 150.9600 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.0800 150.4750 139.2200 150.9600 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.0000 150.4750 140.1400 150.9600 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.4600 150.4750 140.6000 150.9600 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.3800 150.4750 141.5200 150.9600 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.3000 150.4750 142.4400 150.9600 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.7600 150.4750 142.9000 150.9600 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.6800 150.4750 143.8200 150.9600 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.6000 150.4750 144.7400 150.9600 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.0600 150.4750 145.2000 150.9600 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.9800 150.4750 146.1200 150.9600 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.9000 150.4750 147.0400 150.9600 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.3600 150.4750 147.5000 150.9600 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.2800 150.4750 148.4200 150.9600 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.2000 150.4750 149.3400 150.9600 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.1200 150.4750 150.2600 150.9600 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.1200 0.0000 150.2600 0.4850 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.2000 0.0000 149.3400 0.4850 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.8200 0.0000 147.9600 0.4850 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.4400 0.0000 146.5800 0.4850 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.0600 0.0000 145.2000 0.4850 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.6800 0.0000 143.8200 0.4850 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.3000 0.0000 142.4400 0.4850 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.9200 0.0000 141.0600 0.4850 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.5400 0.0000 139.6800 0.4850 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.6200 0.0000 138.7600 0.4850 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.2400 0.0000 137.3800 0.4850 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.8600 0.0000 136.0000 0.4850 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.4800 0.0000 134.6200 0.4850 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.1000 0.0000 133.2400 0.4850 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.7200 0.0000 131.8600 0.4850 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.3400 0.0000 130.4800 0.4850 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.9600 0.0000 129.1000 0.4850 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.0400 0.0000 128.1800 0.4850 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.6600 0.0000 126.8000 0.4850 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.2800 0.0000 125.4200 0.4850 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.9000 0.0000 124.0400 0.4850 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.5200 0.0000 122.6600 0.4850 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.1400 0.0000 121.2800 0.4850 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.7600 0.0000 119.9000 0.4850 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.3800 0.0000 118.5200 0.4850 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.4600 0.0000 117.6000 0.4850 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.0800 0.0000 116.2200 0.4850 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.7000 0.0000 114.8400 0.4850 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.3200 0.0000 113.4600 0.4850 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.9400 0.0000 112.0800 0.4850 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.5600 0.0000 110.7000 0.4850 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.1800 0.0000 109.3200 0.4850 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.8000 0.0000 107.9400 0.4850 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.8800 0.0000 107.0200 0.4850 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.5000 0.0000 105.6400 0.4850 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.1200 0.0000 104.2600 0.4850 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.7400 0.0000 102.8800 0.4850 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.3600 0.0000 101.5000 0.4850 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.5715 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.7495 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.9800 0.0000 100.1200 0.4850 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.7455 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.6195 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 98.6000 0.0000 98.7400 0.4850 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.8099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.9415 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 97.2200 0.0000 97.3600 0.4850 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.3809 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.6785 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 96.3000 0.0000 96.4400 0.4850 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.3165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.3565 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 94.9200 0.0000 95.0600 0.4850 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.9959 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.7535 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 93.5400 0.0000 93.6800 0.4850 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.416 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.851 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.6376 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 159.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 47.7256 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 256.052 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 92.1600 0.0000 92.3000 0.4850 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0994 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.5786 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 185.36 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 77.8797 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 417.477 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 90.7800 0.0000 90.9200 0.4850 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1225 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2585 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 4.78041 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.1047 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 89.4000 0.0000 89.5400 0.4850 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.3238 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.222 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 32.8931 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 159.316 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.498027 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2641 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 33.4879 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 163.443 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.588117 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.7698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 84.576 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 69.0054 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 353.929 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.588117 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 88.0200 0.0000 88.1600 0.4850 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.6533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.8045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 23.9939 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 118.929 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 86.6400 0.0000 86.7800 0.4850 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.1341 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 60.1755 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 100.203 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 487.869 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.7468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.12 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 133.417 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 666.067 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 85.7200 0.0000 85.8600 0.4850 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.97 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.3096 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 14.2108 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 77.9099 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 84.3400 0.0000 84.4800 0.4850 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2702 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.19 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.7356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 180.864 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 75.9811 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 407.351 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 82.9600 0.0000 83.1000 0.4850 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1132 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.229 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.6967 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 94.848 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 39.8574 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 213.622 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 81.5800 0.0000 81.7200 0.4850 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0994 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.6455 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 153.712 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 64.5169 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 346.198 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 80.2000 0.0000 80.3400 0.4850 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3484 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.581 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.265 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.8305 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 144.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 60.4291 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 324.396 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 78.8200 0.0000 78.9600 0.4850 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.6697 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.0795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.0628 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.272 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 111.583 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 585.734 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.9776 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 123.488 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 163.335 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 863.86 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 77.4400 0.0000 77.5800 0.4850 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.4812 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 86.891 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 142.64 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 699.897 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.4229 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.384 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 168.368 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 838.149 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.815487 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.4376 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 88.608 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 205.389 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1037.72 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.815487 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 76.0600 0.0000 76.2000 0.4850 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1132 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.7607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.5573 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 121.712 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 50.8047 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 274.126 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 75.1400 0.0000 75.2800 0.4850 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.1346 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 95.158 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 188.006 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 925.008 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 1.08254 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.4852 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.52 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 382.333 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1968.82 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.4 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.4998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.136 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 403.728 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2083.99 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.4 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 73.7600 0.0000 73.9000 0.4850 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.7961 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.4655 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 101.556 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 503.694 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.31746 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.0188 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.904 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 117.364 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 589.064 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.31746 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 72.3800 0.0000 72.5200 0.4850 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0994 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.775 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.2562 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 211.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 88.4149 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 475.784 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 71.0000 0.0000 71.1400 0.4850 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.1557 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.2835 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 112.347 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 557.806 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.31746 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.4668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.96 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 126.912 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 636.544 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.31746 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 69.6200 0.0000 69.7600 0.4850 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3556 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.617 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.597 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 229.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 346.008 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1820.06 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 5.07937 LAYER via4  ;
    ANTENNADIFFAREA 0.429 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 48.928 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 77.232 LAYER met5  ;
    ANTENNAGATEAREA 0.444 LAYER met5  ;
    ANTENNAMAXAREACAR 456.206 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 1994.01 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 68.2400 0.0000 68.3800 0.4850 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.839 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.3565 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 39.0912 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 210.595 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 66.8600 0.0000 67.0000 0.4850 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.5383 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 117.079 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 186.812 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 929.194 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.31746 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.9848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.056 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 204.796 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1026.17 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.31746 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 65.4800 0.0000 65.6200 0.4850 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.368 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 89.7754 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 435.73 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 101.164 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 500.175 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.6837 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 100.112 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 143.245 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 725.652 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 64.5600 0.0000 64.7000 0.4850 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3484 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.581 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.9824 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 189.987 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 988.806 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.8857 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 175.856 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 264.054 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1384.88 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.22143 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 63.1800 0.0000 63.3200 0.4850 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.4828 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 81.781 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 130.816 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 649.056 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.31746 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.135 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.52 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 139.824 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 700.802 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.634921 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 143.389 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 720.874 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.634921 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 61.8000 0.0000 61.9400 0.4850 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6118 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.898 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.4291 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 90.216 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 72.9614 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 368.189 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 3.11922 LAYER via4  ;
    ANTENNADIFFAREA 0.429 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 12.496 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 22.584 LAYER met5  ;
    ANTENNAGATEAREA 0.444 LAYER met5  ;
    ANTENNAMAXAREACAR 101.106 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 419.054 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 60.4200 0.0000 60.5600 0.4850 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.9216 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.221 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 75.8373 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 366.897 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 77.8286 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 381.246 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.1497 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 145.264 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 138.977 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 708.417 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 59.0400 0.0000 59.1800 0.4850 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.441 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.044 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.2716 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 157.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 65.927 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 353.73 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 57.6600 0.0000 57.8000 0.4850 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.1257 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.3925 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 11.5444 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 57.1903 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 56.2800 0.0000 56.4200 0.4850 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.3633 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.5805 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 14.3318 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 71.1273 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 54.9000 0.0000 55.0400 0.4850 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3249 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.1295 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 30.4295 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 141.815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.498027 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.0868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.6 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 41.8863 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 203.977 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.498027 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 53.9800 0.0000 54.1200 0.4850 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.5455 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 27.9596 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 129.465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.498027 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.3378 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.272 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 35.4771 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 170.618 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.498027 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 52.6000 0.0000 52.7400 0.4850 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.84 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.813 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 86.0595 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 418.008 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 88.0833 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 432.357 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.4708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.856 LAYER met4  ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 115.629 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 550.262 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 6.12222 LAYER via4  ;
    ANTENNADIFFAREA 0.429 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 23.536 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 39.144 LAYER met5  ;
    ANTENNAGATEAREA 1.109 LAYER met5  ;
    ANTENNAMAXAREACAR 136.852 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 585.559 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 51.2200 0.0000 51.3600 0.4850 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.4483 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.1335 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 49.8400 0.0000 49.9800 0.4850 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.9077 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.1345 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.7225 LAYER met2  ;
    ANTENNAMAXAREACAR 5.10843 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.0264 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.0293848 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.4984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.736 LAYER met3  ;
    ANTENNAGATEAREA 9.1575 LAYER met3  ;
    ANTENNAMAXAREACAR 6.03646 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 30.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0293848 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 48.4600 0.0000 48.6000 0.4850 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.9175 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.2325 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.7225 LAYER met2  ;
    ANTENNAMAXAREACAR 18.7228 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 89.118 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.41888 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.4984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.736 LAYER met3  ;
    ANTENNAGATEAREA 9.1575 LAYER met3  ;
    ANTENNAMAXAREACAR 19.6509 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 94.2216 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.41888 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 47.0800 0.0000 47.2200 0.4850 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.8979 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.9875 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.7225 LAYER met2  ;
    ANTENNAMAXAREACAR 5.10483 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.9725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.0293848 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.4984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.736 LAYER met3  ;
    ANTENNAGATEAREA 9.1575 LAYER met3  ;
    ANTENNAMAXAREACAR 6.03286 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 30.076 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0293848 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 45.7000 0.0000 45.8400 0.4850 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.92 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 44.3200 0.0000 44.4600 0.4850 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.018 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 43.4000 0.0000 43.5400 0.4850 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 42.0200 0.0000 42.1600 0.4850 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 40.6400 0.0000 40.7800 0.4850 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4301 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.1405 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 39.2600 0.0000 39.4000 0.4850 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 37.8800 0.0000 38.0200 0.4850 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 36.5000 0.0000 36.6400 0.4850 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 35.1200 0.0000 35.2600 0.4850 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.018 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 33.7400 0.0000 33.8800 0.4850 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.018 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 32.8200 0.0000 32.9600 0.4850 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 31.4400 0.0000 31.5800 0.4850 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 30.0600 0.0000 30.2000 0.4850 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 28.6800 0.0000 28.8200 0.4850 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 27.3000 0.0000 27.4400 0.4850 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 25.9200 0.0000 26.0600 0.4850 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 24.5400 0.0000 24.6800 0.4850 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.018 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 23.1600 0.0000 23.3000 0.4850 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.018 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 22.2400 0.0000 22.3800 0.4850 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 20.8600 0.0000 21.0000 0.4850 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 19.4800 0.0000 19.6200 0.4850 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 18.1000 0.0000 18.2400 0.4850 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 16.7200 0.0000 16.8600 0.4850 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 15.3400 0.0000 15.4800 0.4850 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 13.9600 0.0000 14.1000 0.4850 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.018 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 12.5800 0.0000 12.7200 0.4850 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.018 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 11.6600 0.0000 11.8000 0.4850 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 10.2800 0.0000 10.4200 0.4850 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 8.9000 0.0000 9.0400 0.4850 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 7.5200 0.0000 7.6600 0.4850 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 6.1400 0.0000 6.2800 0.4850 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 4.7600 0.0000 4.9000 0.4850 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.969 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 3.3800 0.0000 3.5200 0.4850 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.018 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2.0000 0.0000 2.1400 0.4850 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3762 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.773 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1.0800 0.0000 1.2200 0.4850 ;
    END
  END io_oeb[0]
  PIN irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3112 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.33 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 148.3400 0.4850 148.4800 ;
    END
  END irq[2]
  PIN irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 149.0200 0.4850 149.1600 ;
    END
  END irq[1]
  PIN irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 150.0400 0.4850 150.1800 ;
    END
  END irq[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.0000 39.8800 0.4800 40.3600 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 45.3200 0.4800 45.8000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 50.7600 0.4800 51.2400 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 56.2000 0.4800 56.6800 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 61.6400 0.4800 62.1200 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 67.0800 0.4800 67.5600 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 72.5200 0.4800 73.0000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 77.9600 0.4800 78.4400 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 83.4000 0.4800 83.8800 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 88.8400 0.4800 89.3200 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 94.2800 0.4800 94.7600 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 99.7200 0.4800 100.2000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 105.1600 0.4800 105.6400 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 110.6000 0.4800 111.0800 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 39.8800 150.8800 40.3600 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 45.3200 150.8800 45.8000 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 50.7600 150.8800 51.2400 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 56.2000 150.8800 56.6800 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 61.6400 150.8800 62.1200 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 67.0800 150.8800 67.5600 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 72.5200 150.8800 73.0000 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 77.9600 150.8800 78.4400 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 83.4000 150.8800 83.8800 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 88.8400 150.8800 89.3200 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 94.2800 150.8800 94.7600 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 99.7200 150.8800 100.2000 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 105.1600 150.8800 105.6400 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 110.6000 150.8800 111.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 40.0200 0.0000 43.3800 3.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 40.0200 147.6000 43.3800 150.9600 ;
    END
    PORT
      LAYER met4 ;
        RECT 67.2200 0.0000 70.5800 3.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 67.2200 147.6000 70.5800 150.9600 ;
    END
    PORT
      LAYER met4 ;
        RECT 94.4200 0.0000 97.7800 3.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 94.4200 147.6000 97.7800 150.9600 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT 40.0200 0.0000 43.3800 150.9600 ;
        RECT 67.2200 0.0000 70.5800 150.9600 ;
        RECT 94.4200 0.0000 97.7800 150.9600 ;
        RECT 39.8550 56.2000 43.3800 56.6800 ;
        RECT 39.8550 39.8800 43.3800 40.3600 ;
        RECT 39.8550 50.7600 43.3800 51.2400 ;
        RECT 39.8550 45.3200 43.3800 45.8000 ;
        RECT 39.8550 72.5200 43.3800 73.0000 ;
        RECT 39.8550 67.0800 43.3800 67.5600 ;
        RECT 39.8550 61.6400 43.3800 62.1200 ;
        RECT 39.8550 94.2800 43.3800 94.7600 ;
        RECT 39.8550 77.9600 43.3800 78.4400 ;
        RECT 39.8550 88.8400 43.3800 89.3200 ;
        RECT 39.8550 83.4000 43.3800 83.8800 ;
        RECT 39.8550 110.6000 43.3800 111.0800 ;
        RECT 39.8550 105.1600 43.3800 105.6400 ;
        RECT 39.8550 99.7200 43.3800 100.2000 ;
    END
# end of P/G power stripe data as pin

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.0000 42.6000 0.4800 43.0800 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 48.0400 0.4800 48.5200 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 53.4800 0.4800 53.9600 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 58.9200 0.4800 59.4000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 64.3600 0.4800 64.8400 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 69.8000 0.4800 70.2800 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 75.2400 0.4800 75.7200 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 80.6800 0.4800 81.1600 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 86.1200 0.4800 86.6000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 91.5600 0.4800 92.0400 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 97.0000 0.4800 97.4800 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 102.4400 0.4800 102.9200 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.0000 107.8800 0.4800 108.3600 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 42.6000 150.8800 43.0800 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 48.0400 150.8800 48.5200 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 53.4800 150.8800 53.9600 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 58.9200 150.8800 59.4000 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 64.3600 150.8800 64.8400 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 69.8000 150.8800 70.2800 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 75.2400 150.8800 75.7200 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 80.6800 150.8800 81.1600 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 86.1200 150.8800 86.6000 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 91.5600 150.8800 92.0400 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 97.0000 150.8800 97.4800 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 102.4400 150.8800 102.9200 ;
    END
    PORT
      LAYER met1 ;
        RECT 150.4000 107.8800 150.8800 108.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.6200 0.0000 56.9800 3.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.6200 147.6000 56.9800 150.9600 ;
    END
    PORT
      LAYER met4 ;
        RECT 80.8200 0.0000 84.1800 3.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 80.8200 147.6000 84.1800 150.9600 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT 53.6200 0.0000 56.9800 150.9600 ;
        RECT 80.8200 0.0000 84.1800 150.9600 ;
    END
# end of P/G power stripe data as pin

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.0000 0.0000 150.8800 150.9600 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 150.8800 150.9600 ;
    LAYER met2 ;
      RECT 0.0000 0.0000 150.8800 150.9600 ;
    LAYER met3 ;
      RECT 0.0000 0.0000 150.8800 150.9600 ;
    LAYER met4 ;
      RECT 0.0000 0.0000 150.8800 150.9600 ;
    LAYER met5 ;
      RECT 0.0000 0.0000 150.8800 150.9600 ;
  END
END user_proj_example

END LIBRARY
