##
## LEF for PtnCells ;
## created by Innovus v17.11-s080_1 on Tue Jun 22 11:43:10 2021
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO user_project_wrapper
  CLASS BLOCK ;
  SIZE 2920.0000 BY 3520.0000 ;
  FOREIGN user_project_wrapper 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 457.553 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2441.69 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.2358 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 97.728 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.492 LAYER met4  ;
    ANTENNAMAXAREACAR 37.0646 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 198.634 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2.7100 -4.8000 3.2700 2.4000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 51.4909 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 257.057 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 121.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 651.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 3.04906 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 19.2201 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 8.2300 -4.8000 8.7900 2.4000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 50.3389 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 251.415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 116.152 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 619.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 110.575 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 544.789 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 26.1700 -4.8000 26.7300 2.4000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 53.1165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 265.303 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 72.436 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 386.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 136.083 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 688.627 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 20.1900 -4.8000 20.7500 2.4000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.2611 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 261.026 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 115.192 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 614.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.504 LAYER met4  ;
    ANTENNAMAXAREACAR 96.4147 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 474.976 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 32.1500 -4.8000 32.7100 2.4000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.815 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.367 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 83.3492 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 408.076 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 126.4500 -4.8000 127.0100 2.4000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 53.0814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 265.118 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3135 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 44.4318 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 221.163 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 102.9900 -4.8000 103.5500 2.4000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 49.3421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 246.432 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.294 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 119.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 101.79 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 522.266 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 79.5300 -4.8000 80.0900 2.4000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.137 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 260.288 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.1588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.4128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.672 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 98.1532 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 506.69 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 55.6100 -4.8000 56.1700 2.4000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9633 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.5375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.2218 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 146.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.944 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 60.0079 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 303.139 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 617.2700 -4.8000 617.8300 2.4000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.4551 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 76.7935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 58.3318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 307.448 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 5.872 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 12.648 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met5  ;
    ANTENNAMAXAREACAR 83.7522 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 344.927 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 599.3300 -4.8000 599.8900 2.4000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0775 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.1085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 43.2888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 231.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.3798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 34.5953 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 176.291 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 581.8500 -4.8000 582.4100 2.4000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 67.9813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 339.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 48.9024 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 243.701 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 563.9100 -4.8000 564.4700 2.4000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0826 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 234.009 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1248.98 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.1604 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 216.808 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 7.44 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 15 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met5  ;
    ANTENNAMAXAREACAR 91.0939 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 355.824 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 546.4300 -4.8000 546.9900 2.4000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3249 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 137.59 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 734.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.6166 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.896 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 42.1424 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 217.626 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 528.4900 -4.8000 529.0500 2.4000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.3927 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.3835 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 43.3986 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 212.388 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 511.0100 -4.8000 511.5700 2.4000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.2735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 62.2708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 333.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.3318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 34.4523 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 175.511 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 493.0700 -4.8000 493.6300 2.4000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.5409 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 77.3605 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 64.0531 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 315.705 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 475.5900 -4.8000 476.1500 2.4000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 38.458 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 207.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.2558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.168 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 29.3164 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 158.255 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 457.6500 -4.8000 458.2100 2.4000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7305 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.4485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3032 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 50.3561 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 260.569 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 439.7100 -4.8000 440.2700 2.4000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.3029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.2355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 61.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 331.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.6614 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.272 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 25.4734 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 135.261 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 422.2300 -4.8000 422.7900 2.4000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.0337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.8895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 68.362 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 365.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 71.0458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 375.256 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 5.488 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 12.072 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met5  ;
    ANTENNAMAXAREACAR 66.9275 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 273.796 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 404.2900 -4.8000 404.8500 2.4000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.1495 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.4685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 85.4548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 456.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.5848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.256 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 34.6861 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 186.893 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 386.8100 -4.8000 387.3700 2.4000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7929 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 61.3528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 328.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.3828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.512 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 25.6394 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 131.188 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 368.8700 -4.8000 369.4300 2.4000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8902 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.172 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 92.0758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 492.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.4868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.4 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 30.2497 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 163.232 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 351.3900 -4.8000 351.9500 2.4000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9267 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 52.609 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 281.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 35.5372 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 180.976 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 333.4500 -4.8000 334.0100 2.4000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1723 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.2285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 77.0218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 407.128 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 11.744 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 25.296 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met5  ;
    ANTENNAMAXAREACAR 86.5614 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 294.905 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 315.9700 -4.8000 316.5300 2.4000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.7932 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 138.215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.7348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 71.6558 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 384.065 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 298.0300 -4.8000 298.5900 2.4000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.1351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.2785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 68.386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 365.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 56.7958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 299.256 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 21.968 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 40.632 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met5  ;
    ANTENNAMAXAREACAR 108.339 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 254.271 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 280.0900 -4.8000 280.6500 2.4000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.1823 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 90.6325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 64.4338 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 344.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 16.5008 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 83.7292 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 262.6100 -4.8000 263.1700 2.4000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.4785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 82.1135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 44.743 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 239.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 88.3271 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 467.083 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 244.6700 -4.8000 245.2300 2.4000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.0735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 184.648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 985.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.6426 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 36.368 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 38.6552 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 205.224 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 227.1900 -4.8000 227.7500 2.4000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7327 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.3845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 41.5006 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 222.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 3.43758 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 20.2343 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.2500 -4.8000 209.8100 2.4000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2887 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.1645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 74.2744 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 393.416 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 9.184 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 17.616 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met5  ;
    ANTENNAMAXAREACAR 112.551 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 459.026 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 191.7700 -4.8000 192.3300 2.4000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.0063 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 84.7525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 64.36 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 343.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 49.5868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 260.808 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 15.984 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 31.656 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met5  ;
    ANTENNAMAXAREACAR 114.53 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 378.913 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 173.8300 -4.8000 174.3900 2.4000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3137 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 194.152 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1035.94 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 40.8236 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 221.657 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 156.3500 -4.8000 156.9100 2.4000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1063 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.2525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 282.561 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1507.93 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.2928 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 66.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 49.6679 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 266.796 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 138.4100 -4.8000 138.9700 2.4000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9227 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.2715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 240.846 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1285.45 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 42.7138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 224.152 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 13.904 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 28.536 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met5  ;
    ANTENNAMAXAREACAR 86.4204 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 262.873 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 114.9500 -4.8000 115.5100 2.4000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5887 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.6645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 310.302 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1655.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.7938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 84.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 63.8133 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 342.238 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 91.0300 -4.8000 91.5900 2.4000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.4847 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 92.1445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.1048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.904 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 137.248 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 209.712 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 201.184 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 307.405 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 67.5700 -4.8000 68.1300 2.4000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9113 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 456.261 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2434.33 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.4388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.144 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 30.0558 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 162.198 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 43.6500 -4.8000 44.2100 2.4000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.4133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 65.9868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 352.4 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 611.2900 -4.8000 611.8500 2.4000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.7095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.2685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 61.21 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 326.92 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.6838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 222.784 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 593.8100 -4.8000 594.3700 2.4000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.6235 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 72.8385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 59.8506 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 320.144 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 575.8700 -4.8000 576.4300 2.4000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7543 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.6105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 283.225 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1511 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 60.7398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 324.416 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 557.9300 -4.8000 558.4900 2.4000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 227.59 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1214.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.45345 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 44.512 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 70.608 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 540.4500 -4.8000 541.0100 2.4000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0325 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 292.853 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1562.35 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 522.5100 -4.8000 523.0700 2.4000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2739 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.0905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 62.518 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 333.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 61.5918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 328.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 505.0300 -4.8000 505.5900 2.4000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0597 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.0195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.42 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.04 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.4608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.928 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 487.0900 -4.8000 487.6500 2.4000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5225 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.3335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 53.368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 285.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 63.8988 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 341.264 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 469.6100 -4.8000 470.1700 2.4000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.3167 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.3045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 64.1928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 342.832 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 451.6700 -4.8000 452.2300 2.4000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.2175 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 77.0208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 411.248 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 434.1900 -4.8000 434.7500 2.4000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.3699 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.5705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 61.69 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 329.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 50.2926 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 269.168 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 416.2500 -4.8000 416.8100 2.4000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.3768 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.4645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 69.6198 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 371.776 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 398.3100 -4.8000 398.8700 2.4000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7509 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.4755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 78.943 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 421.496 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.8838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 293.184 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 380.8300 -4.8000 381.3900 2.4000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.4585 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.0135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 65.2998 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.736 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 362.8900 -4.8000 363.4500 2.4000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.5363 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.4025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.229 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3924 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.776 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 6.976 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 14.304 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 345.4100 -4.8000 345.9700 2.4000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.2423 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.9325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 39.8406 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 213.424 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 327.4700 -4.8000 328.0300 2.4000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.8353 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 164.048 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 309.9900 -4.8000 310.5500 2.4000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.6379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 163.062 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 292.0500 -4.8000 292.6100 2.4000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4522 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.982 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 67.6 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 361 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 62.0928 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 331.632 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 274.5700 -4.8000 275.1300 2.4000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.1857 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.6495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 65.4318 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 349.44 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 256.6300 -4.8000 257.1900 2.4000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.7323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 78.3825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 52.447 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 280.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.6136 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 142.88 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.1500 -4.8000 239.7100 2.4000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.5299 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.4785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 47.6328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 254.512 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 221.2100 -4.8000 221.7700 2.4000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 81.2735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 64.2798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 343.296 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 203.2700 -4.8000 203.8300 2.4000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.2577 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.8915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 65.0178 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 347.232 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 185.7900 -4.8000 186.3500 2.4000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0757 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.9815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 58.978 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 315.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 42.4398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 226.816 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 167.8500 -4.8000 168.4100 2.4000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 282.32 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1507.12 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 150.3700 -4.8000 150.9300 2.4000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4957 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 300.77 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1604.58 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 132.4300 -4.8000 132.9900 2.4000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5945 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 291.754 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1556.49 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.0588 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 176.784 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 108.9700 -4.8000 109.5300 2.4000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5947 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 285.917 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1525.36 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 85.0500 -4.8000 85.6100 2.4000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.3731 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.5865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 172.087 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 918.736 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 61.5900 -4.8000 62.1500 2.4000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3189 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.3305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 219.61 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1171.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 52.9428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 282.832 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 38.1300 -4.8000 38.6900 2.4000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 448.992 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2395.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.536 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 50.5499 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 253.761 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 14.2100 -4.8000 14.7700 2.4000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0396 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.919 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 57.0492 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 306.144 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 623.2500 -4.8000 623.8100 2.4000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0291 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 69.3534 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 371.296 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 605.3100 -4.8000 605.8700 2.4000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8621 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.0315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 65.464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 349.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.1428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 321.232 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 587.8300 -4.8000 588.3900 2.4000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2415 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.9285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 54.8218 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 293.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.4408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 77.488 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 569.8900 -4.8000 570.4500 2.4000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 278.966 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1488.29 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 552.4100 -4.8000 552.9700 2.4000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1427 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.5525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 289.227 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1543.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.6748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 270.736 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 534.4700 -4.8000 535.0300 2.4000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 28.8025 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 143.776 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 516.5300 -4.8000 517.0900 2.4000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.7619 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.5305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 72.3606 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 386.864 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 499.0500 -4.8000 499.6100 2.4000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6079 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.7605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.725 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.45345 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.429 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 78.736 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 121.944 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 481.1100 -4.8000 481.6700 2.4000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.3523 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.1815 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 463.6300 -4.8000 464.1900 2.4000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9797 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 445.6900 -4.8000 446.2500 2.4000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.7715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 48.0048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 256.496 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 428.2100 -4.8000 428.7700 2.4000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7409 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.4255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 53.779 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 287.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.1848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 257.456 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 410.2700 -4.8000 410.8300 2.4000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.6243 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.8425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 392.7900 -4.8000 393.3500 2.4000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.9631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 64.5365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 36.832 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 196.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.9828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.92 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.429 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 58.864 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 92.136 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 374.8500 -4.8000 375.4100 2.4000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.4803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 82.0575 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 357.3700 -4.8000 357.9300 2.4000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.3561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 121.384 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.5958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.648 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 339.4300 -4.8000 339.9900 2.4000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.2131 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 130.721 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 321.4900 -4.8000 322.0500 2.4000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.9159 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 79.1175 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 304.0100 -4.8000 304.5700 2.4000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.4225 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.8335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.1648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 124.016 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 286.0700 -4.8000 286.6300 2.4000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2773 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.7488 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.464 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 268.5900 -4.8000 269.1500 2.4000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.1399 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.3555 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 250.6500 -4.8000 251.2100 2.4000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.2605 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.0235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 57.2028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 305.552 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 233.1700 -4.8000 233.7300 2.4000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8599 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.0205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 79.2486 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 423.6 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 215.2300 -4.8000 215.7900 2.4000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.9011 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.0635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 35.497 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 189.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.024 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.429 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 48.928 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 77.232 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 197.7500 -4.8000 198.3100 2.4000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5721 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.5815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 68.7018 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 366.88 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 179.8100 -4.8000 180.3700 2.4000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.894 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 161.8700 -4.8000 162.4300 2.4000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.2307 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 80.8745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 68.5668 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 366.16 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 144.3900 -4.8000 144.9500 2.4000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.2289 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 85.8655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 34.7568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 185.84 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 120.9300 -4.8000 121.4900 2.4000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7599 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.5205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 254.222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1356.32 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 97.0100 -4.8000 97.5700 2.4000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.1524 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.3075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 148.862 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 794.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.0748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.536 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 73.5500 -4.8000 74.1100 2.4000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.0613 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 80.0275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 37.0548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 198.096 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 49.6300 -4.8000 50.1900 2.4000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2403 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.9225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 235.618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1257.1 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.5058 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 131.168 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2881.3900 -4.8000 2881.9500 2.4000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.0888 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 105.018 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 32.7318 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 175.04 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2863.4500 -4.8000 2864.0100 2.4000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.3801 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 86.6215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.15 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.6746 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.08 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 120.256 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 184.224 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 2845.5100 -4.8000 2846.0700 2.4000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 85.5295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 104.855 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 559.696 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2828.0300 -4.8000 2828.5900 2.4000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2051 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.7465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 236.648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1262.59 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2810.0900 -4.8000 2810.6500 2.4000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.6155 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 102.799 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 77.83 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 415.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.4128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.672 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2792.6100 -4.8000 2793.1700 2.4000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8649 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.0455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 118.618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 633.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 28.3248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 151.536 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2774.6700 -4.8000 2775.2300 2.4000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.3981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 71.7115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 53.9428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 288.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.3618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.608 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 52.048 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 81.912 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 2757.1900 -4.8000 2757.7500 2.4000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0019 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.7305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 124.57 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 664.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.8368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.808 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 43.408 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 68.952 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 2739.2500 -4.8000 2739.8100 2.4000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7215 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.3285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 144.349 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 770.8 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2721.7700 -4.8000 2722.3300 2.4000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.8899 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.1705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 89.3538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 477.024 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2703.8300 -4.8000 2704.3900 2.4000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.2161 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.8015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 104.585 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 558.256 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2685.8900 -4.8000 2686.4500 2.4000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.1631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 95.3435 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2668.4100 -4.8000 2668.9700 2.4000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6519 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.1415 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2650.4700 -4.8000 2651.0300 2.4000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.9871 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 109.421 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.1408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.888 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2632.9900 -4.8000 2633.5500 2.4000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6971 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.2065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 63.8268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 340.88 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2615.0500 -4.8000 2615.6100 2.4000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5679 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6035 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2597.5700 -4.8000 2598.1300 2.4000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9661 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7125 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2579.6300 -4.8000 2580.1900 2.4000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.2267 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 125.78 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2562.1500 -4.8000 2562.7100 2.4000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.3885 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 116.589 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2544.2100 -4.8000 2544.7700 2.4000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.2479 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.004 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2526.7300 -4.8000 2527.2900 2.4000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.8701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 124.072 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.6948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.176 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2508.7900 -4.8000 2509.3500 2.4000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.1529 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 125.486 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.6838 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.784 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2490.8500 -4.8000 2491.4100 2.4000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.0151 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.84 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2473.3700 -4.8000 2473.9300 2.4000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7015 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3895 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2455.4300 -4.8000 2455.9900 2.4000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.2659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 96.0505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.47 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.2688 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 49.904 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2437.9500 -4.8000 2438.5100 2.4000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.5383 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.5735 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2420.0100 -4.8000 2420.5700 2.4000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2325 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0445 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2402.5300 -4.8000 2403.0900 2.4000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.2743 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 111.136 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2384.5900 -4.8000 2385.1500 2.4000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.1259 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 95.3505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.0522 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.16 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2367.1100 -4.8000 2367.6700 2.4000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.3469 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.6065 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2349.1700 -4.8000 2349.7300 2.4000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.2339 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 90.9335 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2331.2300 -4.8000 2331.7900 2.4000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.0457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 114.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2313.7500 -4.8000 2314.3100 2.4000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2501 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.1325 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2295.8100 -4.8000 2296.3700 2.4000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.5763 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 117.646 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2278.3300 -4.8000 2278.8900 2.4000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.8461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.9415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.403 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.0568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 155.44 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2260.3900 -4.8000 2260.9500 2.4000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5893 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.8285 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2242.9100 -4.8000 2243.4700 2.4000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.7263 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.3525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 59.458 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 317.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.048 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 54.448 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 85.512 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 2224.9700 -4.8000 2225.5300 2.4000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.5847 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.6875 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2207.4900 -4.8000 2208.0500 2.4000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0849 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.1885 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2189.5500 -4.8000 2190.1100 2.4000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9709 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.5755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.8238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.072 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 292.912 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 443.208 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 2172.0700 -4.8000 2172.6300 2.4000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.2093 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 85.7675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.172 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.5538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 115.424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2154.1300 -4.8000 2154.6900 2.4000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.9881 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 84.8225 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2136.1900 -4.8000 2136.7500 2.4000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.5217 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.329 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.2608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.528 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2118.7100 -4.8000 2119.2700 2.4000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9643 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.7035 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2100.7700 -4.8000 2101.3300 2.4000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.4673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 111.983 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2083.2900 -4.8000 2083.8500 2.4000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.7467 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 93.3975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.5958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.648 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2065.3500 -4.8000 2065.9100 2.4000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.1939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.7335 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2047.8700 -4.8000 2048.4300 2.4000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.8235 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.9995 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2029.9300 -4.8000 2030.4900 2.4000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 28.4313 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 141.802 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2012.4500 -4.8000 2013.0100 2.4000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.1547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 85.6555 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1994.5100 -4.8000 1995.0700 2.4000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.9287 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 109.365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.9768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 69.68 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1976.5700 -4.8000 1977.1300 2.4000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.7057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 83.2405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.6488 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.264 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1959.0900 -4.8000 1959.6500 2.4000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.2033 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 90.7375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.816 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1941.1500 -4.8000 1941.7100 2.4000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.8051 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 78.9075 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1923.6700 -4.8000 1924.2300 2.4000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.9026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 94.234 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.48 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 120.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.3708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.448 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1905.7300 -4.8000 1906.2900 2.4000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.1677 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 80.7205 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1888.2500 -4.8000 1888.8100 2.4000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.9863 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 89.6525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 86.437 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 461.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.8368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 143.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1870.3100 -4.8000 1870.8700 2.4000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.9651 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 74.7075 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1852.8300 -4.8000 1853.3900 2.4000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.4103 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 76.9335 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1834.8900 -4.8000 1835.4500 2.4000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.7461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 83.5695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 161.122 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 859.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 25.4208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 136.048 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1817.4100 -4.8000 1817.9700 2.4000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8699 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 74.2315 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1799.4700 -4.8000 1800.0300 2.4000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.6428 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 132.699 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.4078 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 34.0113 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 184.352 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1781.5300 -4.8000 1782.0900 2.4000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.4255 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 96.8485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 36.184 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 193.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.5538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 115.424 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.492 LAYER met4  ;
    ANTENNAMAXAREACAR 118.85 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 634.881 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.267073 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1764.0500 -4.8000 1764.6100 2.4000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.3497 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 71.5225 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 137.542 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 683.499 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1746.1100 -4.8000 1746.6700 2.4000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.6197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 92.561 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.619 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 3.91758 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 24.695 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1728.6300 -4.8000 1729.1900 2.4000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.097 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 165.088 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.4851 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 163.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.936 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 5.65576 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 32.0646 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1710.6900 -4.8000 1711.2500 2.4000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.8063 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 88.8055 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 152.611 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 758.845 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1693.2100 -4.8000 1693.7700 2.4000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.2623 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 91.1505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 55.876 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 298.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.1994 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 87.808 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 76.9135 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 411.935 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1675.2700 -4.8000 1675.8300 2.4000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.6435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 102.939 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 32.3506 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 173.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.8238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.072 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 138.352 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 211.368 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 202.803 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 309.833 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 1657.7900 -4.8000 1658.3500 2.4000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.1003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.2225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.543 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.4954 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 287.928 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 21.328 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 35.832 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met5  ;
    ANTENNAMAXAREACAR 86.1737 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 144.776 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 1639.8500 -4.8000 1640.4100 2.4000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.3009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.0425 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 46.6929 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 228.598 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1621.9100 -4.8000 1622.4700 2.4000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.7877 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.593 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.166 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.3008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.616 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 155.248 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 236.712 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 227.57 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 346.983 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 1604.4300 -4.8000 1604.9900 2.4000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.4651 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 77.1645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 88.789 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 474.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 28.0408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 145.896 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 20.736 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 38.784 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met5  ;
    ANTENNAMAXAREACAR 145.653 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 470.388 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 1586.4900 -4.8000 1587.0500 2.4000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.1235 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 75.4565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 57.6976 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 309.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.0118 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 59.2 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 44.4921 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 239.192 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1569.0100 -4.8000 1569.5700 2.4000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0987 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.3325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.723 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 169.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.024 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 413.84 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 628.44 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 629.699 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 1019.93 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 1551.0700 -4.8000 1551.6300 2.4000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3741 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.535 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 115.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.2158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.496 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.4347 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 321.968 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 490.632 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6822 LAYER met5  ;
    ANTENNAMAXAREACAR 487.22 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 776.015 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 1533.5900 -4.8000 1534.1500 2.4000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8893 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.2855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 63.0106 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 337.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2954 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 5.23394 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 33.6162 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1515.6500 -4.8000 1516.2100 2.4000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 145.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3064 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.712 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 85.1188 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 450.461 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1498.1700 -4.8000 1498.7300 2.4000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.3018 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 100.758 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.3518 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.68 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 66.0679 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 354.263 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1480.2300 -4.8000 1480.7900 2.4000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.6456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 167.713 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.0548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.096 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 40.6255 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 218.57 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1462.7500 -4.8000 1463.3100 2.4000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3525 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.35 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 1.95879 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 12.3475 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1444.8100 -4.8000 1445.3700 2.4000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.9867 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 84.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.177 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.5796 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 14.463 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 80.9374 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1426.8700 -4.8000 1427.4300 2.4000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2621 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.0315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.3096 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 40.082 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 213.167 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1409.3900 -4.8000 1409.9500 2.4000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5558 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.382 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.7688 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.904 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 67.7527 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 363.248 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1391.4500 -4.8000 1392.0100 2.4000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.7659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 178.314 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.8348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.256 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 43.777 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 235.378 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1373.9700 -4.8000 1374.5300 2.4000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.0129 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 159.786 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.3506 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.144 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 51.5333 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 271.717 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1356.0300 -4.8000 1356.5900 2.4000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.5251 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 77.3465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.5388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.344 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 50.6618 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 272.097 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1338.5500 -4.8000 1339.1100 2.4000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.2695 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 71.1865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.8658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.7128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 116.272 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 94.0784 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 499.521 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1320.6100 -4.8000 1321.1700 2.4000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.7349 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.3955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.5708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.848 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 60.0489 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 308.651 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1303.1300 -4.8000 1303.6900 2.4000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.8821 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 164.014 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 33.1091 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 164.658 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1285.1900 -4.8000 1285.7500 2.4000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.1805 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 165.624 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.7088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.584 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 63.4291 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 325.737 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1267.2500 -4.8000 1267.8100 2.4000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.4939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 166.978 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.4888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.744 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 34.2982 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 184.824 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1249.7700 -4.8000 1250.3300 2.4000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.0811 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 165.126 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 13.7641 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 66.7535 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1231.8300 -4.8000 1232.3900 2.4000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.8237 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 163.958 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 150.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.7248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.336 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 18.5354 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 93.5394 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1214.3500 -4.8000 1214.9100 2.4000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.0575 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 165.126 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 54.1528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 289.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 1.95879 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 12.3475 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1196.4100 -4.8000 1196.9700 2.4000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.7895 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 168.829 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1178.9300 -4.8000 1179.4900 2.4000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.2283 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 165.98 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 43.7238 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 233.664 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1160.9900 -4.8000 1161.5500 2.4000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.6579 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 168.172 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1143.5100 -4.8000 1144.0700 2.4000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 30.6801 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.283 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1125.5700 -4.8000 1126.1300 2.4000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.1677 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 170.678 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 59.6358 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 318.528 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1107.6300 -4.8000 1108.1900 2.4000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.7429 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 173.596 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1090.1500 -4.8000 1090.7100 2.4000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.8261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 168.969 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 71.4558 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 381.568 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1072.2100 -4.8000 1072.7700 2.4000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.4055 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 171.91 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1054.7300 -4.8000 1055.2900 2.4000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.9485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 174.507 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1036.7900 -4.8000 1037.3500 2.4000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.3901 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 171.672 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.9448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 128.176 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1019.3100 -4.8000 1019.8700 2.4000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.458 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 172.011 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 45.7368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 244.4 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1001.3700 -4.8000 1001.9300 2.4000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.3817 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 171.79 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 983.8900 -4.8000 984.4500 2.4000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.5717 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 177.74 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 965.9500 -4.8000 966.5100 2.4000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.2021 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 175.732 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.4988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.464 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 948.4700 -4.8000 949.0300 2.4000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.0215 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 174.99 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 930.5300 -4.8000 931.0900 2.4000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.7149 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 173.456 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 912.5900 -4.8000 913.1500 2.4000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.4527 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 177.146 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 895.1100 -4.8000 895.6700 2.4000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.4205 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 176.824 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 53.3028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 284.752 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 877.1700 -4.8000 877.7300 2.4000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.4289 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 177.026 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 859.6900 -4.8000 860.2500 2.4000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.3365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 176.404 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.3328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.912 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 841.7500 -4.8000 842.3100 2.4000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 38.3003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 191.383 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 824.2700 -4.8000 824.8300 2.4000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.9525 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 179.645 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 806.3300 -4.8000 806.8900 2.4000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 36.2381 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 181.072 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 788.8500 -4.8000 789.4100 2.4000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.8615 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 179.029 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.0368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 770.9100 -4.8000 771.4700 2.4000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.6687 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 173.064 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.0468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 112.72 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 752.9700 -4.8000 753.5300 2.4000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 30.1829 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 150.678 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 735.4900 -4.8000 736.0500 2.4000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.7789 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 178.616 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.7948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 143.376 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 717.5500 -4.8000 718.1100 2.4000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 36.2059 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 180.751 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.5438 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 152.704 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 700.0700 -4.8000 700.6300 2.4000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.1071 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 155.418 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 682.1300 -4.8000 682.6900 2.4000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 36.8051 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 183.746 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.1228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.792 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 664.6500 -4.8000 665.2100 2.4000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.3171 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 171.188 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.7548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.496 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 646.7100 -4.8000 647.2700 2.4000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 37.0737 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 185.132 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 629.2300 -4.8000 629.7900 2.4000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4055 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 71.6835 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2886.9100 -4.8000 2887.4700 2.4000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.5175 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.3085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 241.292 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1287.36 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2869.4300 -4.8000 2869.9900 2.4000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.0503 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 134.908 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2851.4900 -4.8000 2852.0500 2.4000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.1197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.3195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 79.8148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 426.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2834.0100 -4.8000 2834.5700 2.4000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.3065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.2925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 118.108 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 630.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.5898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 275.616 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2816.0700 -4.8000 2816.6300 2.4000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 51.0879 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 255.16 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 47.893 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 255.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.3118 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 156.8 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2798.5900 -4.8000 2799.1500 2.4000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 49.0394 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 244.853 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2780.6500 -4.8000 2781.2100 2.4000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 53.6919 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 268.18 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 64.9788 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 347.024 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2763.1700 -4.8000 2763.7300 2.4000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 51.2069 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 255.756 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 39.2628 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 209.872 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2745.2300 -4.8000 2745.7900 2.4000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 71.9881 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 359.426 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.7778 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.952 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2727.2900 -4.8000 2727.8500 2.4000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.2039 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 170.74 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 57.025 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 304.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.8986 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 208.4 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2709.8100 -4.8000 2710.3700 2.4000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.0839 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 95.1405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 75.1428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 401.232 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2691.8700 -4.8000 2692.4300 2.4000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.3583 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 236.512 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 66.49 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 355.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.1508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.608 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2674.3900 -4.8000 2674.9500 2.4000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.9771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 64.6065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 105.598 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 563.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.9448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 288.176 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2656.4500 -4.8000 2657.0100 2.4000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.1341 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.3915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 67.858 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 362.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.7518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 164.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2638.9700 -4.8000 2639.5300 2.4000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8169 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.9135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 314.092 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1676.1 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2621.0300 -4.8000 2621.5900 2.4000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6291 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.9745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 48.493 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 259.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 79.2558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 423.168 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2603.5500 -4.8000 2604.1100 2.4000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 38.8323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.882 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.7128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.272 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2585.6100 -4.8000 2586.1700 2.4000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 38.6741 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 193.092 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.184 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2567.6700 -4.8000 2568.2300 2.4000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 41.7487 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 208.282 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2550.1900 -4.8000 2550.7500 2.4000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.1529 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 195.486 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.6988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.864 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2532.2500 -4.8000 2532.8100 2.4000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.692 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.762 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.6938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.504 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2514.7700 -4.8000 2515.3300 2.4000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.3266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 216.118 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.5158 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.888 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2496.8300 -4.8000 2497.3900 2.4000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.5591 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.5165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.026 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 68.9508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 368.208 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2479.3500 -4.8000 2479.9100 2.4000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.4519 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.0335 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2461.4100 -4.8000 2461.9700 2.4000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.0937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.1245 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2443.9300 -4.8000 2444.4900 2.4000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 51.2393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 255.734 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2425.9900 -4.8000 2426.5500 2.4000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.7099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 113.271 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.8168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 202.16 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2408.5100 -4.8000 2409.0700 2.4000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.7609 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 223.29 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.6368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2390.5700 -4.8000 2391.1300 2.4000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.0352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 214.543 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.0628 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.472 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2372.6300 -4.8000 2373.1900 2.4000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.8541 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.9265 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2355.1500 -4.8000 2355.7100 2.4000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 40.3863 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 201.652 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.0188 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.904 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2337.2100 -4.8000 2337.7700 2.4000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.6871 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.0915 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2319.7300 -4.8000 2320.2900 2.4000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.8273 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.9105 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2301.7900 -4.8000 2302.3500 2.4000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.6633 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.9725 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2284.3100 -4.8000 2284.8700 2.4000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 41.5243 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 207.225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.6948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.176 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2266.3700 -4.8000 2266.9300 2.4000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.7521 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.4815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 64.291 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 343.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 65.1558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 347.968 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2248.8900 -4.8000 2249.4500 2.4000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.0895 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2230.9500 -4.8000 2231.5100 2.4000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.0239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.8405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 69.052 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 368.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 70.0806 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 374.704 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2213.0100 -4.8000 2213.5700 2.4000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.3647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 226.544 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.727 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.7598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.856 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2195.5300 -4.8000 2196.0900 2.4000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.5263 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.4055 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2177.5900 -4.8000 2178.1500 2.4000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.2613 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.9625 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2160.1100 -4.8000 2160.6700 2.4000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.3949 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.6955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.4688 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.304 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2142.1700 -4.8000 2142.7300 2.4000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8579 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 84.0105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.2128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 284.272 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2124.6900 -4.8000 2125.2500 2.4000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8475 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.0015 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2106.7500 -4.8000 2107.3100 2.4000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.8881 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.9785 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2089.2700 -4.8000 2089.8300 2.4000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.0013 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.7275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.335 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.92 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 65.9118 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 352 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2071.3300 -4.8000 2071.8900 2.4000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.5481 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.4615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 94.351 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 503.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 69.4206 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 371.184 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2053.8500 -4.8000 2054.4100 2.4000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 27.6262 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.669 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2035.9100 -4.8000 2036.4700 2.4000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.5689 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 72.5445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.59 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 126.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 61.5516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 329.216 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2017.9700 -4.8000 2018.5300 2.4000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.4712 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 77.077 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.805 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.8548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 79.696 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2000.4900 -4.8000 2001.0500 2.4000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.1731 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.576 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.9198 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 117.376 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1982.5500 -4.8000 1983.1100 2.4000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 51.5163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 257.302 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 74.2476 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 396.928 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1965.0700 -4.8000 1965.6300 2.4000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.3081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 96.3795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 159.832 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 852.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.024 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.336 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 201.616 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 306.264 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 1947.1300 -4.8000 1947.6900 2.4000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 51.7487 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 258.465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 90.1176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.568 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1929.6500 -4.8000 1930.2100 2.4000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.4937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 87.3075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 91.522 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 488.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.5636 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.488 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.336 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 94.864 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 146.136 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 1911.7100 -4.8000 1912.2700 2.4000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.4553 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 217.116 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 125.083 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 667.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.2788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 61.832 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.336 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 162.64 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 247.8 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 1894.2300 -4.8000 1894.7900 2.4000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 43.8713 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 219.012 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1876.2900 -4.8000 1876.8500 2.4000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.3091 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 81.2665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.751 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.2998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.736 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1858.3500 -4.8000 1858.9100 2.4000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.2413 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 60.9805 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1840.8700 -4.8000 1841.4300 2.4000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.7946 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 83.629 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1822.9300 -4.8000 1823.4900 2.4000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.6405 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 262.923 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 79.8798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 426.496 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1805.4500 -4.8000 1806.0100 2.4000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 85.5295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.45345 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.336 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 38.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 62.328 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 1787.5100 -4.8000 1788.0700 2.4000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 47.3454 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 236.383 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1770.0300 -4.8000 1770.5900 2.4000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.0025 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 239.852 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 134.708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 718.912 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1752.0900 -4.8000 1752.6500 2.4000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.3441 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 241.56 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 75.4158 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 402.688 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1734.6100 -4.8000 1735.1700 2.4000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.6647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 243.162 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 130.946 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 699.792 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1716.6700 -4.8000 1717.2300 2.4000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.9089 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.2655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.4308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.768 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1699.1900 -4.8000 1699.7500 2.4000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.8317 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 238.997 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 71.971 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 384.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1681.2500 -4.8000 1681.8100 2.4000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 73.8 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 368.774 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1663.3100 -4.8000 1663.8700 2.4000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.1547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 260.495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 61.2948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 327.376 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1645.8300 -4.8000 1646.3900 2.4000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 69.0582 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 345.065 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1627.8900 -4.8000 1628.4500 2.4000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 49.7959 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 248.818 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 90.7278 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 484.352 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1610.4100 -4.8000 1610.9700 2.4000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.0173 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 229.926 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 77.077 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 411.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.7788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.624 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1592.4700 -4.8000 1593.0300 2.4000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 57.7155 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 288.298 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.7648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.216 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1574.9900 -4.8000 1575.5500 2.4000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.8533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 263.988 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.1588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.984 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1557.0500 -4.8000 1557.6100 2.4000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.7119 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 228.281 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 58.7886 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 314.48 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1539.5700 -4.8000 1540.1300 2.4000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.9947 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 229.694 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.7296 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.832 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1521.6300 -4.8000 1522.1900 2.4000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.0635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 230.156 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 70.1518 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 375.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.2098 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.256 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1503.6900 -4.8000 1504.2500 2.4000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.9113 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 224.396 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.354 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.1656 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.824 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1486.2100 -4.8000 1486.7700 2.4000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.2698 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 96.005 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1468.2700 -4.8000 1468.8300 2.4000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.3315 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.4965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.405 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.8688 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 245.104 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1450.7900 -4.8000 1451.3500 2.4000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 28.0103 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 139.772 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.5028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.152 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1432.8500 -4.8000 1433.4100 2.4000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.1383 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.5305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.402 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 67.3596 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 360.192 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1415.3700 -4.8000 1415.9300 2.4000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.5325 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.2655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.251 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.1598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.656 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1397.4300 -4.8000 1397.9900 2.4000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 24.636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 122.836 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1379.9500 -4.8000 1380.5100 2.4000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 38.4792 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 192.052 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1362.0100 -4.8000 1362.5700 2.4000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 28.5604 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 142.576 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1344.0700 -4.8000 1344.6300 2.4000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 30.7494 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 153.167 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1326.5900 -4.8000 1327.1500 2.4000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.2353 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 145.898 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.0188 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.904 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1308.6500 -4.8000 1309.2100 2.4000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 46.2956 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 231.252 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1291.1700 -4.8000 1291.7300 2.4000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.6133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 237.906 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.6418 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.56 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1273.2300 -4.8000 1273.7900 2.4000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 46.0826 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 230.069 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1255.7500 -4.8000 1256.3100 2.4000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.1087 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 225.382 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.0818 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 150.24 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1237.8100 -4.8000 1238.3700 2.4000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 52.6276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 262.794 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1220.3300 -4.8000 1220.8900 2.4000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 53.5992 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 267.652 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1202.3900 -4.8000 1202.9500 2.4000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.9849 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 229.646 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.0168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.56 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met3  ;
    ANTENNAMAXAREACAR 50.6543 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 245.362 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.472349 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1184.9100 -4.8000 1185.4700 2.4000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.5075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 227.258 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.407 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 141.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.1786 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 252.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 54.3219 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 290.248 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1166.9700 -4.8000 1167.5300 2.4000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.0404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 230.041 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 52.5108 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 280.528 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 101.765 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 522.807 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.461485 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1149.0300 -4.8000 1149.5900 2.4000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.4157 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 221.918 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 58.816 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 314.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.1564 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 172.432 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 78.2347 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 411.372 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1131.5500 -4.8000 1132.1100 2.4000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 49.0536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 244.517 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met2  ;
    ANTENNAMAXAREACAR 90.3025 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 440.227 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.715332 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.339 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.608 LAYER met3  ;
    ANTENNAGATEAREA 0.621 LAYER met3  ;
    ANTENNAMAXAREACAR 102.12 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 504.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.779744 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.0107 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.856 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 115.522 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 576.105 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.779744 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1113.6100 -4.8000 1114.1700 2.4000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 56.9915 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 284.399 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.896 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 6.39893 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 36.0054 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.0535475 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.4258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.408 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 13.6624 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 75.3735 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0535475 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1096.1300 -4.8000 1096.6900 2.4000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.2089 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 75.8835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.3538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 45.024 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 96.0721 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 486.678 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.778944 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1078.1900 -4.8000 1078.7500 2.4000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.5455 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 242.449 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.1946 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 136.52 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.429 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 25.744 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 42.456 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.441 LAYER met5  ;
    ANTENNAMAXAREACAR 58.3764 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 96.2721 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 1060.7100 -4.8000 1061.2700 2.4000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 50.3795 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 251.618 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.947 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.5994 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 180.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 38.6867 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 207.954 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1042.7700 -4.8000 1043.3300 2.4000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.0003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 229.722 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.2147 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 25.7225 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 137.81 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1025.2900 -4.8000 1025.8500 2.4000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.6113 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 227.896 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 56.4988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 302.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.9233 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 123.664 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 88.4383 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 462.298 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.638219 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1007.3500 -4.8000 1007.9100 2.4000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.0573 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 235.008 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 54.6778 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 292.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.2668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.56 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 7.0506 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 38.2329 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 989.4100 -4.8000 989.9700 2.4000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 232.666 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.613 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.5842 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 175.184 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 57.9684 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 300.498 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 971.9300 -4.8000 972.4900 2.4000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.4937 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 242.189 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.2115 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 178.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 44.4598 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 238.372 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 953.9900 -4.8000 954.5500 2.4000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 61.4924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 306.894 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.8732 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.256 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met3  ;
    ANTENNAMAXAREACAR 14.9555 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 80.6999 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.0402212 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.5478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.392 LAYER met4  ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 21.5395 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 116.288 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0402212 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 936.5100 -4.8000 937.0700 2.4000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.5621 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 227.532 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.1726 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.528 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 94.6286 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 467.194 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.41387 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 918.5700 -4.8000 919.1300 2.4000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.2339 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 236.008 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 116.856 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 624.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.0034 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 219.616 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 41.2302 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 220.831 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 901.0900 -4.8000 901.6500 2.4000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.6495 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 237.968 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.97 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.192 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 84.9096 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 441.16 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.665585 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 883.1500 -4.8000 883.7100 2.4000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.8679 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 239.061 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 57.0718 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 305.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.8687 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 138.432 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 26.0118 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 139.198 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 865.6700 -4.8000 866.2300 2.4000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 56.1305 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 280.255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.5941 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.6144 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 228.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 57.0474 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 306.142 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 847.7300 -4.8000 848.2900 2.4000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 50.5643 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 252.542 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.7949 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 93.6103 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 502.921 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.31746 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.2078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.912 LAYER met4  ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 106.891 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 574.225 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.31746 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 830.2500 -4.8000 830.8100 2.4000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 53.1135 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 265.171 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.747 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.2035 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 19.0141 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 102.661 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 812.3100 -4.8000 812.8700 2.4000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 53.9031 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 269.118 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.402 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.7186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 95.44 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 17.8166 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 95.9678 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 794.3700 -4.8000 794.9300 2.4000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 38.1461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 190.334 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.8895 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 117.68 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 29.3032 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 157.537 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 776.8900 -4.8000 777.4500 2.4000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.5145 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 227.294 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.024 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.429 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 118.816 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 182.064 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met5  ;
    ANTENNAMAXAREACAR 173.276 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 439.93 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 758.9500 -4.8000 759.5100 2.4000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 40.0363 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 199.902 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.1618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 108 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 26.9904 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 144.578 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 741.4700 -4.8000 742.0300 2.4000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.4669 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 227.056 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.1382 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 151.952 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 28.2938 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 152.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 723.5300 -4.8000 724.0900 2.4000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 66.135 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 329.987 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.57 LAYER met2  ;
    ANTENNAMAXAREACAR 122.994 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 604.543 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 706.0500 -4.8000 706.6100 2.4000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.4311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 236.876 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 62.2488 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 332.464 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met3  ;
    ANTENNAMAXAREACAR 89.8685 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 459.938 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.626729 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 688.1100 -4.8000 688.6700 2.4000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.3475 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 231.458 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 32.8798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 176.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.7828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 95.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 23.8056 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 127.593 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 670.6300 -4.8000 671.1900 2.4000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.9305 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 244.374 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.1836 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 151.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.9017 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 90.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8175 LAYER met4  ;
    ANTENNAMAXAREACAR 20.6749 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 110.835 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 652.6900 -4.8000 653.2500 2.4000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 53.0605 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 265.023 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.1736 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 151.2 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1325 LAYER met4  ;
    ANTENNAMAXAREACAR 24.8774 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 133.51 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 634.7500 -4.8000 635.3100 2.4000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 62.8703 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 314.233 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2892.8900 -4.8000 2893.4500 2.4000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 54.0293 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 270.029 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2875.4100 -4.8000 2875.9700 2.4000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 37.1369 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 185.406 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 32.1348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 171.856 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2857.4700 -4.8000 2858.0300 2.4000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.4137 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 226.951 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2839.9900 -4.8000 2840.5500 2.4000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 49.1377 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 245.41 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 73.7436 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 394.24 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2822.0500 -4.8000 2822.6100 2.4000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.8599 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 234.02 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.7628 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 169.872 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2804.1100 -4.8000 2804.6700 2.4000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.6533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 242.988 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 35.932 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 192.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.9748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.336 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2786.6300 -4.8000 2787.1900 2.4000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 49.1489 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 245.465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 101.081 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 539.568 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2768.6900 -4.8000 2769.2500 2.4000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.5476 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 242.459 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 59.0868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 315.6 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2751.2100 -4.8000 2751.7700 2.4000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.8499 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 233.852 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.8768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2733.2700 -4.8000 2733.8300 2.4000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.0437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 230.1 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2715.7900 -4.8000 2716.3500 2.4000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 60.2943 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 301.354 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2697.8500 -4.8000 2698.4100 2.4000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 60.8599 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 304.021 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2680.3700 -4.8000 2680.9300 2.4000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 61.7377 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 308.57 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2662.4300 -4.8000 2662.9900 2.4000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 60.4315 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 302.039 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2644.9500 -4.8000 2645.5100 2.4000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 61.1931 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 305.847 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2627.0100 -4.8000 2627.5700 2.4000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.3957 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 241.7 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.457 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 130.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.8216 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.656 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2609.0700 -4.8000 2609.6300 2.4000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 42.7439 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 213.44 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.2288 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.232 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 108.544 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 166.656 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 2591.5900 -4.8000 2592.1500 2.4000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.3003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 226.222 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.5348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 168.656 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2573.6500 -4.8000 2574.2100 2.4000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.6843 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 223.303 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2556.1700 -4.8000 2556.7300 2.4000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 49.5297 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 247.37 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 33.7908 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 180.688 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2538.2300 -4.8000 2538.7900 2.4000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 49.1419 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 245.43 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 124.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2520.7500 -4.8000 2521.3100 2.4000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.7169 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 218.306 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.8808 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.168 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2502.8100 -4.8000 2503.3700 2.4000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 58.6703 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 293.233 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2485.3300 -4.8000 2485.8900 2.4000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 59.3423 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 296.594 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2467.3900 -4.8000 2467.9500 2.4000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.6993 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 228.378 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2449.4500 -4.8000 2450.0100 2.4000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 225.69 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2431.9700 -4.8000 2432.5300 2.4000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.9499 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 229.632 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2414.0300 -4.8000 2414.5900 2.4000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.4801 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 222.24 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 291.487 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1555.06 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.9968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.12 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2396.5500 -4.8000 2397.1100 2.4000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.9381 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 219.572 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2378.6100 -4.8000 2379.1700 2.4000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.5523 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 227.482 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.1048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.904 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 71.008 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 110.352 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 2361.1300 -4.8000 2361.6900 2.4000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.3437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 226.439 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.865 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.1018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.68 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2343.1900 -4.8000 2343.7500 2.4000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 58.1971 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 290.867 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2325.7100 -4.8000 2326.2700 2.4000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 59.7511 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 298.638 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2307.7700 -4.8000 2308.3300 2.4000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 55.4391 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 277.078 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2290.2900 -4.8000 2290.8500 2.4000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 54.1357 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 270.561 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2272.3500 -4.8000 2272.9100 2.4000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 56.1139 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 280.451 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2254.4100 -4.8000 2254.9700 2.4000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 57.1191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 285.478 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2236.9300 -4.8000 2237.4900 2.4000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 57.6903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 288.333 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2218.9900 -4.8000 2219.5500 2.4000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 56.5479 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 282.621 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2201.5100 -4.8000 2202.0700 2.4000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 58.7375 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 293.57 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2183.5700 -4.8000 2184.1300 2.4000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 58.3763 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 291.763 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2166.0900 -4.8000 2166.6500 2.4000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 55.7863 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 278.814 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2148.1500 -4.8000 2148.7100 2.4000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 55.1059 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 275.411 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2130.6700 -4.8000 2131.2300 2.4000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.5443 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.4425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 68.1528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 363.952 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2112.7300 -4.8000 2113.2900 2.4000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.4713 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 222.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2094.7900 -4.8000 2095.3500 2.4000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.8289 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 218.866 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.771 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.2418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 50.968 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 121.792 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 186.528 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 2077.3100 -4.8000 2077.8700 2.4000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.4441 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 222.092 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2059.3700 -4.8000 2059.9300 2.4000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.6527 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 232.984 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 36.5928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 195.632 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2041.8900 -4.8000 2042.4500 2.4000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.9787 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 234.658 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2023.9500 -4.8000 2024.5100 2.4000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.9163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 229.302 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 36.046 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 192.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.4128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.672 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2006.4700 -4.8000 2007.0300 2.4000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.7003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 163.383 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1988.5300 -4.8000 1989.0900 2.4000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 50.7685 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 253.606 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1971.0500 -4.8000 1971.6100 2.4000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 54.6551 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 273.158 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1953.1100 -4.8000 1953.6700 2.4000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 50.9465 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 254.615 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1935.6300 -4.8000 1936.1900 2.4000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.1869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 235.742 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.1248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.136 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1917.6900 -4.8000 1918.2500 2.4000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.9935 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 244.85 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1899.7500 -4.8000 1900.3100 2.4000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 51.9307 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 259.535 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1882.2700 -4.8000 1882.8300 2.4000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 51.5443 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 257.604 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1864.3300 -4.8000 1864.8900 2.4000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 54.2559 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 271.043 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1846.8500 -4.8000 1847.4100 2.4000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.2613 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 235.952 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1828.9100 -4.8000 1829.4700 2.4000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0826 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.2065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 75.2424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 402.704 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1811.4300 -4.8000 1811.9900 2.4000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.9605 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 234.406 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.278 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.0074 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 118.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met4  ;
    ANTENNAMAXAREACAR 83.4333 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 446.761 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.413208 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1793.4900 -4.8000 1794.0500 2.4000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.1919 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 235.798 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 98.815 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 527.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.315 LAYER met4  ;
    ANTENNAMAXAREACAR 36.7717 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 185.485 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.417143 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1776.0100 -4.8000 1776.5700 2.4000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.4653 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 232.165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 99.826 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 532.872 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 22.2014 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 113.026 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265454 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1758.0700 -4.8000 1758.6300 2.4000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.4901 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 237.29 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 83.911 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 447.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 28.2019 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 144.465 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265454 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1740.1300 -4.8000 1740.6900 2.4000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.9901 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 234.672 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.2156 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.424 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 8.1 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 41.4313 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1722.6500 -4.8000 1723.2100 2.4000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 49.4513 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 246.978 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2739 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.856 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 17.3831 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 85.5394 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1704.7100 -4.8000 1705.2700 2.4000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.0979 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 235.21 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 13.4837 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 66.8747 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1687.2300 -4.8000 1687.7900 2.4000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 51.1019 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 255.23 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.0598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.456 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 10.2218 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 55.4667 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1669.2900 -4.8000 1669.8500 2.4000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 50.3641 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 251.542 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.2228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 2.4703 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 14.1253 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1651.8100 -4.8000 1652.3700 2.4000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.7694 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.621 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 42.5153 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 210.936 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1633.8700 -4.8000 1634.4300 2.4000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.1853 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 260.53 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.9276 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.888 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 17.6584 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 89.1313 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1616.3900 -4.8000 1616.9500 2.4000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 53.3431 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 266.318 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 19.6256 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 97.4484 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1598.4500 -4.8000 1599.0100 2.4000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.5679 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 242.561 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.4778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 72.352 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 27.2279 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 146.166 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1580.9700 -4.8000 1581.5300 2.4000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.1923 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 240.447 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6828 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.112 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 18.4024 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 91.8929 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1563.0300 -4.8000 1563.5900 2.4000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.5807 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 222.624 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.3516 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 162.816 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 76.6414 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 403.881 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1545.0900 -4.8000 1545.6500 2.4000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.5703 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 197.69 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.6 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.0684 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 65.776 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 40.6956 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 215.547 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265454 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1527.6100 -4.8000 1528.1700 2.4000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.3087 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 226.264 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.7304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.64 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 35.8987 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 191.945 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1509.6700 -4.8000 1510.2300 2.4000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.5931 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 227.804 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.452 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 9.44576 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 50.2869 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265454 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1492.1900 -4.8000 1492.7500 2.4000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.1365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 225.404 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 13.9369 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 68.8828 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1474.2500 -4.8000 1474.8100 2.4000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.1132 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 145.222 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 59.6024 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 295.997 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1456.7700 -4.8000 1457.3300 2.4000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.6918 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 108.115 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 44.3788 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 220.015 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1438.8300 -4.8000 1439.3900 2.4000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.8812 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 104.062 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 42.7412 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 211.827 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1421.3500 -4.8000 1421.9100 2.4000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.7832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 138.572 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 56.6846 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 281.544 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1403.4100 -4.8000 1403.9700 2.4000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.0908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 110.11 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 45.1848 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 224.045 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1385.4700 -4.8000 1386.0300 2.4000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.821 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.761 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 42.7204 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 211.587 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1367.9900 -4.8000 1368.5500 2.4000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.7709 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 83.4575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 63.7972 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 338.008 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 11.744 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 25.296 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met5  ;
    ANTENNAMAXAREACAR 61.4244 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 238.06 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 1350.0500 -4.8000 1350.6100 2.4000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.7064 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 83.188 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 37.0723 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 183.346 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1332.5700 -4.8000 1333.1300 2.4000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.849 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 138.901 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 56.8176 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 282.209 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1314.6300 -4.8000 1315.1900 2.4000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.0208 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 144.76 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 59.9361 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 297.666 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1297.1500 -4.8000 1297.7100 2.4000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.7429 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 228.553 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.329 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 124.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.5198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 45.7398 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 238.186 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265454 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1279.2100 -4.8000 1279.7700 2.4000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.8573 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 199.126 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.7634 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.816 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 52.0052 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 271.359 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265454 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1261.7300 -4.8000 1262.2900 2.4000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.7723 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 228.701 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 52.234 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 279.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.3258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 28.0246 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 144.408 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265454 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1243.7900 -4.8000 1244.3500 2.4000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.6967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 228.322 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.7408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 159.088 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 78.1653 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 409.798 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1225.8500 -4.8000 1226.4100 2.4000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.5231 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 242.337 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 15.6713 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 77.4384 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.184646 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1208.3700 -4.8000 1208.9300 2.4000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 49.5045 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 247.404 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1190.4300 -4.8000 1190.9900 2.4000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 49.7383 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 248.574 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1172.9500 -4.8000 1173.5100 2.4000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.0153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 234.798 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 39.523 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 211.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1155.0100 -4.8000 1155.5700 2.4000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.1015 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 260.389 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1137.5300 -4.8000 1138.0900 2.4000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 51.2587 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 256.176 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1119.5900 -4.8000 1120.1500 2.4000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 50.0211 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 249.988 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1102.1100 -4.8000 1102.6700 2.4000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.7835 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 243.799 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1084.1700 -4.8000 1084.7300 2.4000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 50.0687 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 250.226 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1066.6900 -4.8000 1067.2500 2.4000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 51.8033 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 258.898 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1048.7500 -4.8000 1049.3100 2.4000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.0989 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 225.334 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 65.941 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 352.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.7388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.952 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 363.712 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 549.408 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 1030.8100 -4.8000 1031.3700 2.4000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.6211 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 227.944 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 49.7796 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 266.432 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1013.3300 -4.8000 1013.8900 2.4000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.0989 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 225.334 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 51.9078 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 277.312 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 995.3900 -4.8000 995.9500 2.4000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.9529 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 229.604 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 78.4356 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 419.264 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 977.9100 -4.8000 978.4700 2.4000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.8465 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 229.072 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 38.7108 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 206.928 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 959.9700 -4.8000 960.5300 2.4000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.3799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 231.738 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 151.73 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 809.696 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 942.4900 -4.8000 943.0500 2.4000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 51.9195 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 259.318 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.041 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 107.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.1358 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.528 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 924.5500 -4.8000 925.1100 2.4000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.0257 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 259.892 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 907.0700 -4.8000 907.6300 2.4000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 50.4915 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 252.34 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 889.1300 -4.8000 889.6900 2.4000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 51.4659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 257.212 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 871.1900 -4.8000 871.7500 2.4000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 51.5779 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 257.611 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.8868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.2 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 853.7100 -4.8000 854.2700 2.4000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.1749 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 235.757 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 835.7700 -4.8000 836.3300 2.4000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.5035 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 242.238 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 49.3368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 263.6 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 818.2900 -4.8000 818.8500 2.4000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 51.6213 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 257.828 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 47.686 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 254.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.45345 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 30.16 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 49.08 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 800.3500 -4.8000 800.9100 2.4000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 54.1509 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 270.358 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.4048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.296 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 782.8700 -4.8000 783.4300 2.4000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.6491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 328.009 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 764.9300 -4.8000 765.4900 2.4000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 53.3069 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 266.255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 65.2548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.496 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 747.4500 -4.8000 748.0100 2.4000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 50.7477 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 253.46 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 65.3448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 348.976 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 729.5100 -4.8000 730.0700 2.4000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.6347 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 262.776 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.9658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.288 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 712.0300 -4.8000 712.5900 2.4000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 50.0029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 249.736 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 42.649 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 227.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.024 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 171.376 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 260.904 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 694.0900 -4.8000 694.6500 2.4000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 60.1163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 300.345 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 676.1500 -4.8000 676.7100 2.4000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.3663 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 241.552 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 37.453 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 200.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 658.6700 -4.8000 659.2300 2.4000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.1885 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 240.663 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.029 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 155.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3924 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.776 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 69.904 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 108.696 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 640.7300 -4.8000 641.2900 2.4000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 62.8212 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 335.512 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 161.5800 2.4000 162.7800 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.5864 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.456 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 357.4200 2.4000 358.6200 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.336 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 552.5800 2.4000 553.7800 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.736 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 813.7000 2.4000 814.9000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.0684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.36 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1074.1400 2.4000 1075.3400 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.304 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1335.2600 2.4000 1336.4600 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 82.5222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 440.584 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1595.7000 2.4000 1596.9000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.0264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 112.136 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1856.1400 2.4000 1857.3400 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2117.2600 2.4000 2118.4600 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.5054 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2377.7000 2.4000 2378.9000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.5392 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 350.008 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2638.8200 2.4000 2640.0200 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 63.7362 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 340.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2899.2600 2.4000 2900.4600 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 81.8622 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 437.064 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 3159.7000 2.4000 3160.9000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 65.6712 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 350.712 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 3420.8200 2.4000 3422.0200 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 475.05 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2374.97 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 51.3138 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 274.144 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 202.3500 3517.6000 202.9100 3524.8000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 475.004 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2374.74 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 61.2468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 327.12 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 527.1100 3517.6000 527.6700 3524.8000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 476.31 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2381.27 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 61.9398 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 330.816 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 851.4100 3517.6000 851.9700 3524.8000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 473.317 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2366.42 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 69.5298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 371.296 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1175.7100 3517.6000 1176.2700 3524.8000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 213.074 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1065.25 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1500.4700 3517.6000 1501.0300 3524.8000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 471.097 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2355.32 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 113.833 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 607.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.7398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1824.7700 3517.6000 1825.3300 3524.8000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 471.274 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2356.09 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.374 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2149.0700 3517.6000 2149.6300 3524.8000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 596.566 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2982.55 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.2428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.432 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2473.8300 3517.6000 2474.3900 3524.8000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 474.246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2370.95 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.2588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 167.184 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2798.1300 3517.6000 2798.6900 3524.8000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 3352.8200 2924.8000 3354.0200 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.3538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 189.024 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 3086.9400 2924.8000 3088.1400 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.848 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2821.0600 2924.8000 2822.2600 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2555.8600 2924.8000 2557.0600 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2289.9800 2924.8000 2291.1800 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2716 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 373.256 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1991.17 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2024.1000 2924.8000 2025.3000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.5076 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.648 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1758.9000 2924.8000 1760.1000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2866 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 325.724 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1737.66 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1493.0200 2924.8000 1494.2200 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 37.4052 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 199.96 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1227.1400 2924.8000 1228.3400 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.0988 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 59.664 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1027.9000 2924.8000 1029.1000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3054 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.624 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 828.6600 2924.8000 829.8600 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.6938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.504 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 629.4200 2924.8000 630.6200 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.2204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 430.1800 2924.8000 431.3800 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 230.9400 2924.8000 232.1400 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.1272 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 177.144 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 32.3800 2924.8000 33.5800 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 363.616 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1939.75 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 96.3000 2.4000 97.5000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.8434 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 111.16 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 292.1400 2.4000 293.3400 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.00165 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.008 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 487.3000 2.4000 488.5000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 30.6634 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 164 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.1766 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.216 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 748.4200 2.4000 749.6200 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.2894 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1008.8600 2.4000 1010.0600 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 63.2532 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 337.816 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1269.9800 2.4000 1271.1800 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 61.5762 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 328.872 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.621 LAYER met3  ;
    ANTENNAMAXAREACAR 142.753 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 746.343 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0644122 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1530.4200 2.4000 1531.6200 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 78.4792 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 419.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.1786 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 252.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 54.3219 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 290.248 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1791.5400 2.4000 1792.7400 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 357.943 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1788.57 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0535475 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2051.9800 2.4000 2053.1800 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.1854 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.3816 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 40.6715 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 217.531 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2312.4200 2.4000 2313.6200 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.7508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 171.016 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.429 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 217.744 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 330.456 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met5  ;
    ANTENNAMAXAREACAR 307.089 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 521.296 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2573.5400 2.4000 2574.7400 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.78735 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.4258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.408 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 7.26345 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 39.3681 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2833.9800 2.4000 2835.1800 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.7458 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.384 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 13.0466 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 71.4645 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 3095.1000 2.4000 3096.3000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.2394 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.12 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.441 LAYER met3  ;
    ANTENNAMAXAREACAR 63.2777 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 311.385 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.94932 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3924 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.776 LAYER met4  ;
    ANTENNAGATEAREA 0.441 LAYER met4  ;
    ANTENNAMAXAREACAR 66.4351 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 319.948 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 2.40057 LAYER via4  ;
    ANTENNADIFFAREA 0.429 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 25.744 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 42.456 LAYER met5  ;
    ANTENNAGATEAREA 0.441 LAYER met5  ;
    ANTENNAMAXAREACAR 124.812 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 416.22 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 3355.5400 2.4000 3356.7400 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 284.632 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1422.88 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.9351 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.5994 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 180.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8685 LAYER met4  ;
    ANTENNAMAXAREACAR 38.6867 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 207.954 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 121.3900 3517.6000 121.9500 3524.8000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 265.521 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1327.43 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.6215 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.584 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 240.619 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1198.52 LAYER met3  ;
    ANTENNAMAXCUTCAR 1.53889 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 445.6900 3517.6000 446.2500 3524.8000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 471.31 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2356.27 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.619 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.6293 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 138.096 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 25.7711 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 138.86 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 770.4500 3517.6000 771.0100 3524.8000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 472.719 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2363.43 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 95.8726 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 512.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 252.267 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1291.42 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.41387 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.2668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.56 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 259.318 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1329.65 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.41387 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1094.7500 3517.6000 1095.3100 3524.8000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 317.879 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1589.12 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.718 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.0014 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 166.272 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 31.1729 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 167.192 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1419.0500 3517.6000 1419.6100 3524.8000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 470.328 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2351.48 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 108.884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 581.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.2115 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 178.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 44.4598 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 238.372 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1743.8100 3517.6000 1744.3700 3524.8000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 476.024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2379.72 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.1372 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.064 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met3  ;
    ANTENNAMAXAREACAR 100.965 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 499.387 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.40054 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.5478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.392 LAYER met4  ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 107.549 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 534.975 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.40054 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 2068.1100 3517.6000 2068.6700 3524.8000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 472.41 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2361.77 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 50.7303 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 271.968 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 103.138 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 538.12 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.346262 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 2392.4100 3517.6000 2392.9700 3524.8000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 288.297 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1441.09 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.0034 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 219.616 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 41.2302 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 220.831 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2717.1700 3517.6000 2717.7300 3524.8000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.3458 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 75.8151 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 389.222 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.3488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 151.664 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 113.765 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 592.253 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.36032 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 3418.7800 2924.8000 3419.9800 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.4294 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.152 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 119.069 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 597.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.8687 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 138.432 LAYER met4  ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 145.081 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 737.15 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 3153.5800 2924.8000 3154.7800 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.6144 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 228.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 57.0474 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 306.142 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2887.7000 2924.8000 2888.9000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.0589 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.176 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 272.363 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1386.83 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.2078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.912 LAYER met4  ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 285.644 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1458.14 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2621.8200 2924.8000 2623.0200 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0857 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.9493 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 145.136 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 127.403 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 651.204 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.99524 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2356.6200 2924.8000 2357.8200 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 392.828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2096.5 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 893.129 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 4709.44 LAYER met4  ;
    ANTENNAMAXCUTCAR 2.17381 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2090.7400 2924.8000 2091.9400 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.5772 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.344 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 262.6 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1359.4 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.8895 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 117.68 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 291.904 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1516.94 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.67778 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1824.8600 2924.8000 1826.0600 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1146 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 310.423 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1656.53 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 353.685 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1877.09 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0804424 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1559.6600 2924.8000 1560.8600 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 40.6962 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 217.96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 95.7831 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 487.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.800698 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.1618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 108 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 122.773 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 631.738 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.800698 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1293.7800 2924.8000 1294.9800 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.0904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 208.944 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.4556 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 104.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met4  ;
    ANTENNAMAXAREACAR 67.3905 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 345.779 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.609043 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1094.5400 2924.8000 1095.7400 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 49.3632 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 263.736 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.57 LAYER met3  ;
    ANTENNAMAXAREACAR 110.183 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 579.319 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0701754 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 895.3000 2924.8000 896.5000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.2484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.32 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9945 LAYER met3  ;
    ANTENNAMAXAREACAR 94.6386 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 473.275 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0402212 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 696.0600 2924.8000 697.2600 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.2014 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.536 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.747 LAYER met3  ;
    ANTENNAMAXAREACAR 78.9031 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 386.604 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.800698 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.7828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 95.312 LAYER met4  ;
    ANTENNAGATEAREA 0.747 LAYER met4  ;
    ANTENNAMAXAREACAR 102.709 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 514.197 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.800698 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 496.8200 2924.8000 498.0200 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.2553 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 135.152 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.57 LAYER met3  ;
    ANTENNAMAXAREACAR 241.3 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1211.57 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.31145 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.9017 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 90.608 LAYER met4  ;
    ANTENNAGATEAREA 0.8175 LAYER met4  ;
    ANTENNAMAXAREACAR 261.975 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1322.4 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.31145 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 297.5800 2924.8000 298.7800 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.1736 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 151.2 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1325 LAYER met4  ;
    ANTENNAMAXAREACAR 24.8774 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 133.51 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 98.3400 2924.8000 99.5400 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2754 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 31.7000 2.4000 32.9000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.0854 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 8.7885 LAYER met4  ;
    ANTENNAMAXAREACAR 4.49378 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 22.8375 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0091028 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 226.8600 2.4000 228.0600 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 8.7885 LAYER met3  ;
    ANTENNAMAXAREACAR 20.4089 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 99.2716 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.348591 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 422.7000 2.4000 423.9000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.1744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 8.7885 LAYER met3  ;
    ANTENNAMAXAREACAR 12.6629 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 63.4667 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0045514 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 683.1400 2.4000 684.3400 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.8094 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 116.312 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 943.5800 2.4000 944.7800 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.2144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.472 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1204.7000 2.4000 1205.9000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7854 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1465.1400 2.4000 1466.3400 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.1774 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.608 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1726.2600 2.4000 1727.4600 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.6274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.008 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1986.7000 2.4000 1987.9000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2247.1400 2.4000 2248.3400 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.256 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2508.2600 2.4000 2509.4600 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 37.6992 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 201.528 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2768.7000 2.4000 2769.9000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.105 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.496 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 3029.8200 2.4000 3031.0200 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.622 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 142.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.1538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.624 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 3290.2600 2.4000 3291.4600 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 301.433 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1507.04 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 40.4300 3517.6000 40.9900 3524.8000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 471.032 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2354.76 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.555 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 364.7300 3517.6000 365.2900 3524.8000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 472.255 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2361 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.409 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 130.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 689.0300 3517.6000 689.5900 3524.8000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 485.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2427.93 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1013.7900 3517.6000 1014.3500 3524.8000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 443.085 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2215.27 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.592 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.0078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 320.512 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1338.0900 3517.6000 1338.6500 3524.8000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 474.513 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2372.4 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 64.729 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 345.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.9644 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.888 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1662.3900 3517.6000 1662.9500 3524.8000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 464.642 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2322.93 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.0748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.9618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1987.1500 3517.6000 1987.7100 3524.8000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 491.83 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2458.9 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2311.4500 3517.6000 2312.0100 3524.8000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 470.877 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2354.1 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.7716 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 181.056 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2635.7500 3517.6000 2636.3100 3524.8000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 59.8182 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 319.496 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 3485.4200 2924.8000 3486.6200 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.088 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 3219.5400 2924.8000 3220.7400 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.2878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.88 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.3365 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 210.112 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 319.008 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2954.3400 2924.8000 2955.5400 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9234 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.5226 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.728 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2688.4600 2924.8000 2689.6600 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9234 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.8978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.8 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.3365 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 167.728 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 255.432 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2422.5800 2924.8000 2423.7800 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2654 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 362.744 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1936.05 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2157.3800 2924.8000 2158.5800 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.8448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.976 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1891.5000 2924.8000 1892.7000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.0228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.592 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1625.6200 2924.8000 1626.8200 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0492 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.728 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1360.4200 2924.8000 1361.6200 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.8244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1161.1800 2924.8000 1162.3800 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 77.4312 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 413.432 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 961.9400 2924.8000 963.1400 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.0124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.728 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 762.7000 2924.8000 763.9000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.4388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.144 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 563.4600 2924.8000 564.6600 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.352 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 364.2200 2924.8000 365.4200 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.337 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.0226 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.728 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 164.9800 2924.8000 166.1800 ;
    END
  END io_oeb[0]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 617.8600 2.4000 619.0600 ;
    END
  END analog_io[28]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 878.9800 2.4000 880.1800 ;
    END
  END analog_io[27]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1139.4200 2.4000 1140.6200 ;
    END
  END analog_io[26]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1399.8600 2.4000 1401.0600 ;
    END
  END analog_io[25]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1660.9800 2.4000 1662.1800 ;
    END
  END analog_io[24]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1921.4200 2.4000 1922.6200 ;
    END
  END analog_io[23]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2182.5400 2.4000 2183.7400 ;
    END
  END analog_io[22]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2442.9800 2.4000 2444.1800 ;
    END
  END analog_io[21]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2703.4200 2.4000 2704.6200 ;
    END
  END analog_io[20]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2964.5400 2.4000 2965.7400 ;
    END
  END analog_io[19]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 3224.9800 2.4000 3226.1800 ;
    END
  END analog_io[18]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 3486.1000 2.4000 3487.3000 ;
    END
  END analog_io[17]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.7700 3517.6000 284.3300 3524.8000 ;
    END
  END analog_io[16]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.0700 3517.6000 608.6300 3524.8000 ;
    END
  END analog_io[15]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.3700 3517.6000 932.9300 3524.8000 ;
    END
  END analog_io[14]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.1300 3517.6000 1257.6900 3524.8000 ;
    END
  END analog_io[13]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.4300 3517.6000 1581.9900 3524.8000 ;
    END
  END analog_io[12]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.7300 3517.6000 1906.2900 3524.8000 ;
    END
  END analog_io[11]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.4900 3517.6000 2231.0500 3524.8000 ;
    END
  END analog_io[10]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.7900 3517.6000 2555.3500 3524.8000 ;
    END
  END analog_io[9]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.0900 3517.6000 2879.6500 3524.8000 ;
    END
  END analog_io[8]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 3286.1800 2924.8000 3287.3800 ;
    END
  END analog_io[7]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 3020.3000 2924.8000 3021.5000 ;
    END
  END analog_io[6]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2755.1000 2924.8000 2756.3000 ;
    END
  END analog_io[5]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2489.2200 2924.8000 2490.4200 ;
    END
  END analog_io[4]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2223.3400 2924.8000 2224.5400 ;
    END
  END analog_io[3]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1958.1400 2924.8000 1959.3400 ;
    END
  END analog_io[2]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1692.2600 2924.8000 1693.4600 ;
    END
  END analog_io[1]
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1426.3800 2924.8000 1427.5800 ;
    END
  END analog_io[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.8700 -4.8000 2899.4300 2.4000 ;
    END
  END user_clock2
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 49.2147 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 245.794 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.675 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 137.4 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2916.8100 -4.8000 2917.3700 2.4000 ;
    END
  END user_irq[2]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.0415 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 239.928 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.299 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.336 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.3124 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 77.744 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2910.8300 -4.8000 2911.3900 2.4000 ;
    END
  END user_irq[1]
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 49.7733 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 248.588 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.336 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 77.9898 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 416.416 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2904.8500 -4.8000 2905.4100 2.4000 ;
    END
  END user_irq[0]
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 2917.6000 158.3800 2962.5000 161.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 158.3800 2.4000 161.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 338.3800 2962.5000 341.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 338.3800 2.4000 341.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 518.3800 2962.5000 521.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 518.3800 2.4000 521.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 698.3800 2962.5000 701.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 698.3800 2.4000 701.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 878.3800 2962.5000 881.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 878.3800 2.4000 881.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1058.3800 2962.5000 1061.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1058.3800 2.4000 1061.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1238.3800 2962.5000 1241.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1238.3800 2.4000 1241.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1418.3800 2962.5000 1421.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1418.3800 2.4000 1421.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1598.3800 2962.5000 1601.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1598.3800 2.4000 1601.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1778.3800 2962.5000 1781.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1778.3800 2.4000 1781.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1958.3800 2962.5000 1961.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1958.3800 2.4000 1961.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2138.3800 2962.5000 2141.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2138.3800 2.4000 2141.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2318.3800 2962.5000 2321.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2318.3800 2.4000 2321.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2498.3800 2962.5000 2501.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2498.3800 2.4000 2501.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2678.3800 2962.5000 2681.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2678.3800 2.4000 2681.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2858.3800 2962.5000 2861.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2858.3800 2.4000 2861.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3038.3800 2962.5000 3041.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 3038.3800 2.4000 3041.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3218.3800 2962.5000 3221.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 3218.3800 2.4000 3221.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3398.3800 2962.5000 3401.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 3398.3800 2.4000 3401.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 3554.2000 2962.5000 3557.2000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2962.5000 -37.5200 2962.5000 -34.5200 ;
    END
    PORT
      LAYER met4 ;
        RECT 153.0200 -37.5200 156.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 153.0200 3517.6000 156.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 333.0200 -37.5200 336.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 333.0200 3517.6000 336.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 513.0200 -37.5200 516.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 513.0200 3517.6000 516.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.0200 -37.5200 696.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.0200 3517.6000 696.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 873.0200 -37.5200 876.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 873.0200 3517.6000 876.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.0200 -37.5200 1056.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.0200 3517.6000 1056.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1233.0200 -37.5200 1236.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1233.0200 3517.6000 1236.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1413.0200 -37.5200 1416.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1413.0200 3517.6000 1416.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1593.0200 -37.5200 1596.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1593.0200 3517.6000 1596.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1773.0200 -37.5200 1776.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1773.0200 3517.6000 1776.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1953.0200 -37.5200 1956.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1953.0200 3517.6000 1956.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2133.0200 -37.5200 2136.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2133.0200 3517.6000 2136.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2313.0200 -37.5200 2316.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2313.0200 3517.6000 2316.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2493.0200 -37.5200 2496.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2493.0200 3517.6000 2496.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2673.0200 -37.5200 2676.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2673.0200 3517.6000 2676.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2853.0200 -37.5200 2856.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2853.0200 3517.6000 2856.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT -42.8800 3557.2000 -39.8800 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2959.5000 -37.5200 2962.5000 3557.2000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT -42.8800 -37.5200 -39.8800 3557.2000 ;
        RECT 2959.5000 -37.5200 2962.5000 3557.2000 ;
      LAYER met5 ;
        RECT -42.8800 -37.5200 2962.5000 -34.5200 ;
        RECT -42.8800 3554.2000 2962.5000 3557.2000 ;
        RECT -42.8800 -37.5300 -39.8800 -34.5100 ;
        RECT 153.0200 -37.5300 156.0200 -34.5100 ;
        RECT 333.0200 -37.5300 336.0200 -34.5100 ;
        RECT 513.0200 -37.5300 516.0200 -34.5100 ;
        RECT 693.0200 -37.5300 696.0200 -34.5100 ;
        RECT 873.0200 -37.5300 876.0200 -34.5100 ;
        RECT 1053.0200 -37.5300 1056.0200 -34.5100 ;
        RECT 1233.0200 -37.5300 1236.0200 -34.5100 ;
        RECT 1413.0200 -37.5300 1416.0200 -34.5100 ;
        RECT 1593.0200 -37.5300 1596.0200 -34.5100 ;
        RECT 1773.0200 -37.5300 1776.0200 -34.5100 ;
        RECT 1953.0200 -37.5300 1956.0200 -34.5100 ;
        RECT 2133.0200 -37.5300 2136.0200 -34.5100 ;
        RECT 2313.0200 -37.5300 2316.0200 -34.5100 ;
        RECT 2493.0200 -37.5300 2496.0200 -34.5100 ;
        RECT 2673.0200 -37.5300 2676.0200 -34.5100 ;
        RECT 2853.0200 -37.5300 2856.0200 -34.5100 ;
        RECT 2959.5000 -37.5300 2962.5000 -34.5100 ;
        RECT -42.8800 878.3700 -39.8800 881.3900 ;
        RECT -42.8800 158.3700 -39.8800 161.3900 ;
        RECT -42.8800 338.3700 -39.8800 341.3900 ;
        RECT -42.8800 518.3700 -39.8800 521.3900 ;
        RECT -42.8800 698.3700 -39.8800 701.3900 ;
        RECT -42.8800 1058.3700 -39.8800 1061.3900 ;
        RECT -42.8800 1238.3700 -39.8800 1241.3900 ;
        RECT -42.8800 1418.3700 -39.8800 1421.3900 ;
        RECT -42.8800 1598.3700 -39.8800 1601.3900 ;
        RECT 2959.5000 878.3700 2962.5000 881.3900 ;
        RECT 2959.5000 158.3700 2962.5000 161.3900 ;
        RECT 2959.5000 338.3700 2962.5000 341.3900 ;
        RECT 2959.5000 518.3700 2962.5000 521.3900 ;
        RECT 2959.5000 698.3700 2962.5000 701.3900 ;
        RECT 2959.5000 1058.3700 2962.5000 1061.3900 ;
        RECT 2959.5000 1238.3700 2962.5000 1241.3900 ;
        RECT 2959.5000 1418.3700 2962.5000 1421.3900 ;
        RECT 2959.5000 1598.3700 2962.5000 1601.3900 ;
        RECT -42.8800 1778.3700 -39.8800 1781.3900 ;
        RECT -42.8800 1958.3700 -39.8800 1961.3900 ;
        RECT -42.8800 2138.3700 -39.8800 2141.3900 ;
        RECT -42.8800 2318.3700 -39.8800 2321.3900 ;
        RECT -42.8800 2498.3700 -39.8800 2501.3900 ;
        RECT -42.8800 2858.3700 -39.8800 2861.3900 ;
        RECT -42.8800 2678.3700 -39.8800 2681.3900 ;
        RECT -42.8800 3038.3700 -39.8800 3041.3900 ;
        RECT -42.8800 3218.3700 -39.8800 3221.3900 ;
        RECT -42.8800 3398.3700 -39.8800 3401.3900 ;
        RECT 2959.5000 1778.3700 2962.5000 1781.3900 ;
        RECT 2959.5000 1958.3700 2962.5000 1961.3900 ;
        RECT 2959.5000 2138.3700 2962.5000 2141.3900 ;
        RECT 2959.5000 2318.3700 2962.5000 2321.3900 ;
        RECT 2959.5000 2498.3700 2962.5000 2501.3900 ;
        RECT 2959.5000 2858.3700 2962.5000 2861.3900 ;
        RECT 2959.5000 2678.3700 2962.5000 2681.3900 ;
        RECT 2959.5000 3038.3700 2962.5000 3041.3900 ;
        RECT 2959.5000 3218.3700 2962.5000 3221.3900 ;
        RECT 2959.5000 3398.3700 2962.5000 3401.3900 ;
        RECT -42.8800 3554.1900 -39.8800 3557.2100 ;
        RECT 153.0200 3554.1900 156.0200 3557.2100 ;
        RECT 333.0200 3554.1900 336.0200 3557.2100 ;
        RECT 513.0200 3554.1900 516.0200 3557.2100 ;
        RECT 693.0200 3554.1900 696.0200 3557.2100 ;
        RECT 873.0200 3554.1900 876.0200 3557.2100 ;
        RECT 1053.0200 3554.1900 1056.0200 3557.2100 ;
        RECT 1233.0200 3554.1900 1236.0200 3557.2100 ;
        RECT 1413.0200 3554.1900 1416.0200 3557.2100 ;
        RECT 1593.0200 3554.1900 1596.0200 3557.2100 ;
        RECT 1773.0200 3554.1900 1776.0200 3557.2100 ;
        RECT 1953.0200 3554.1900 1956.0200 3557.2100 ;
        RECT 2133.0200 3554.1900 2136.0200 3557.2100 ;
        RECT 2313.0200 3554.1900 2316.0200 3557.2100 ;
        RECT 2493.0200 3554.1900 2496.0200 3557.2100 ;
        RECT 2673.0200 3554.1900 2676.0200 3557.2100 ;
        RECT 2853.0200 3554.1900 2856.0200 3557.2100 ;
        RECT 2959.5000 3554.1900 2962.5000 3557.2100 ;
    END
# end of P/G power stripe data as pin

  END vssa2
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 2917.6000 140.3800 2953.1000 143.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 140.3800 2.4000 143.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 320.3800 2953.1000 323.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 320.3800 2.4000 323.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 500.3800 2953.1000 503.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 500.3800 2.4000 503.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 680.3800 2953.1000 683.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 680.3800 2.4000 683.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 860.3800 2953.1000 863.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 860.3800 2.4000 863.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1040.3800 2953.1000 1043.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1040.3800 2.4000 1043.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1220.3800 2953.1000 1223.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1220.3800 2.4000 1223.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1400.3800 2953.1000 1403.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1400.3800 2.4000 1403.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1580.3800 2953.1000 1583.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1580.3800 2.4000 1583.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1760.3800 2953.1000 1763.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1760.3800 2.4000 1763.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1940.3800 2953.1000 1943.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1940.3800 2.4000 1943.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2120.3800 2953.1000 2123.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2120.3800 2.4000 2123.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2300.3800 2953.1000 2303.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2300.3800 2.4000 2303.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2480.3800 2953.1000 2483.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2480.3800 2.4000 2483.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2660.3800 2953.1000 2663.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2660.3800 2.4000 2663.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2840.3800 2953.1000 2843.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2840.3800 2.4000 2843.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3020.3800 2953.1000 3023.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 3020.3800 2.4000 3023.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3200.3800 2953.1000 3203.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 3200.3800 2.4000 3203.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3380.3800 2953.1000 3383.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 3380.3800 2.4000 3383.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 3544.8000 2953.1000 3547.8000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2953.1000 -28.1200 2953.1000 -25.1200 ;
    END
    PORT
      LAYER met4 ;
        RECT 135.0200 -28.1200 138.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 135.0200 3517.6000 138.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 315.0200 -28.1200 318.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 315.0200 3517.6000 318.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 495.0200 -28.1200 498.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 495.0200 3517.6000 498.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.0200 -28.1200 678.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.0200 3517.6000 678.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 855.0200 -28.1200 858.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 855.0200 3517.6000 858.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1035.0200 -28.1200 1038.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1035.0200 3517.6000 1038.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1215.0200 -28.1200 1218.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1215.0200 3517.6000 1218.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1395.0200 -28.1200 1398.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1395.0200 3517.6000 1398.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1575.0200 -28.1200 1578.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1575.0200 3517.6000 1578.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1755.0200 -28.1200 1758.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1755.0200 3517.6000 1758.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1935.0200 -28.1200 1938.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1935.0200 3517.6000 1938.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2115.0200 -28.1200 2118.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2115.0200 3517.6000 2118.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2295.0200 -28.1200 2298.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2295.0200 3517.6000 2298.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2475.0200 -28.1200 2478.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2475.0200 3517.6000 2478.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2655.0200 -28.1200 2658.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2655.0200 3517.6000 2658.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2835.0200 -28.1200 2838.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2835.0200 3517.6000 2838.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT -33.4800 3547.8000 -30.4800 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2950.1000 -28.1200 2953.1000 3547.8000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT -33.4800 -28.1200 -30.4800 3547.8000 ;
        RECT 2950.1000 -28.1200 2953.1000 3547.8000 ;
      LAYER met5 ;
        RECT -33.4800 -28.1200 2953.1000 -25.1200 ;
        RECT -33.4800 3544.8000 2953.1000 3547.8000 ;
        RECT -33.4800 -28.1300 -30.4800 -25.1100 ;
        RECT 135.0200 -28.1300 138.0200 -25.1100 ;
        RECT 315.0200 -28.1300 318.0200 -25.1100 ;
        RECT 495.0200 -28.1300 498.0200 -25.1100 ;
        RECT 675.0200 -28.1300 678.0200 -25.1100 ;
        RECT 855.0200 -28.1300 858.0200 -25.1100 ;
        RECT 1035.0200 -28.1300 1038.0200 -25.1100 ;
        RECT 1395.0200 -28.1300 1398.0200 -25.1100 ;
        RECT 1215.0200 -28.1300 1218.0200 -25.1100 ;
        RECT 1575.0200 -28.1300 1578.0200 -25.1100 ;
        RECT 1755.0200 -28.1300 1758.0200 -25.1100 ;
        RECT 1935.0200 -28.1300 1938.0200 -25.1100 ;
        RECT 2295.0200 -28.1300 2298.0200 -25.1100 ;
        RECT 2115.0200 -28.1300 2118.0200 -25.1100 ;
        RECT 2475.0200 -28.1300 2478.0200 -25.1100 ;
        RECT 2655.0200 -28.1300 2658.0200 -25.1100 ;
        RECT 2835.0200 -28.1300 2838.0200 -25.1100 ;
        RECT 2950.1000 -28.1300 2953.1000 -25.1100 ;
        RECT -33.4800 140.3700 -30.4800 143.3900 ;
        RECT -33.4800 320.3700 -30.4800 323.3900 ;
        RECT -33.4800 500.3700 -30.4800 503.3900 ;
        RECT -33.4800 680.3700 -30.4800 683.3900 ;
        RECT -33.4800 860.3700 -30.4800 863.3900 ;
        RECT -33.4800 1040.3700 -30.4800 1043.3900 ;
        RECT -33.4800 1220.3700 -30.4800 1223.3900 ;
        RECT -33.4800 1400.3700 -30.4800 1403.3900 ;
        RECT -33.4800 1580.3700 -30.4800 1583.3900 ;
        RECT 2950.1000 140.3700 2953.1000 143.3900 ;
        RECT 2950.1000 320.3700 2953.1000 323.3900 ;
        RECT 2950.1000 500.3700 2953.1000 503.3900 ;
        RECT 2950.1000 680.3700 2953.1000 683.3900 ;
        RECT 2950.1000 860.3700 2953.1000 863.3900 ;
        RECT 2950.1000 1040.3700 2953.1000 1043.3900 ;
        RECT 2950.1000 1220.3700 2953.1000 1223.3900 ;
        RECT 2950.1000 1400.3700 2953.1000 1403.3900 ;
        RECT 2950.1000 1580.3700 2953.1000 1583.3900 ;
        RECT -33.4800 1760.3700 -30.4800 1763.3900 ;
        RECT -33.4800 1940.3700 -30.4800 1943.3900 ;
        RECT -33.4800 2120.3700 -30.4800 2123.3900 ;
        RECT -33.4800 2300.3700 -30.4800 2303.3900 ;
        RECT -33.4800 2480.3700 -30.4800 2483.3900 ;
        RECT -33.4800 2660.3700 -30.4800 2663.3900 ;
        RECT -33.4800 2840.3700 -30.4800 2843.3900 ;
        RECT -33.4800 3020.3700 -30.4800 3023.3900 ;
        RECT -33.4800 3200.3700 -30.4800 3203.3900 ;
        RECT -33.4800 3380.3700 -30.4800 3383.3900 ;
        RECT 2950.1000 1760.3700 2953.1000 1763.3900 ;
        RECT 2950.1000 1940.3700 2953.1000 1943.3900 ;
        RECT 2950.1000 2120.3700 2953.1000 2123.3900 ;
        RECT 2950.1000 2300.3700 2953.1000 2303.3900 ;
        RECT 2950.1000 2480.3700 2953.1000 2483.3900 ;
        RECT 2950.1000 2660.3700 2953.1000 2663.3900 ;
        RECT 2950.1000 2840.3700 2953.1000 2843.3900 ;
        RECT 2950.1000 3020.3700 2953.1000 3023.3900 ;
        RECT 2950.1000 3200.3700 2953.1000 3203.3900 ;
        RECT 2950.1000 3380.3700 2953.1000 3383.3900 ;
        RECT -33.4800 3544.7900 -30.4800 3547.8100 ;
        RECT 135.0200 3544.7900 138.0200 3547.8100 ;
        RECT 315.0200 3544.7900 318.0200 3547.8100 ;
        RECT 495.0200 3544.7900 498.0200 3547.8100 ;
        RECT 675.0200 3544.7900 678.0200 3547.8100 ;
        RECT 855.0200 3544.7900 858.0200 3547.8100 ;
        RECT 1035.0200 3544.7900 1038.0200 3547.8100 ;
        RECT 1395.0200 3544.7900 1398.0200 3547.8100 ;
        RECT 1215.0200 3544.7900 1218.0200 3547.8100 ;
        RECT 1575.0200 3544.7900 1578.0200 3547.8100 ;
        RECT 1755.0200 3544.7900 1758.0200 3547.8100 ;
        RECT 1935.0200 3544.7900 1938.0200 3547.8100 ;
        RECT 2295.0200 3544.7900 2298.0200 3547.8100 ;
        RECT 2115.0200 3544.7900 2118.0200 3547.8100 ;
        RECT 2475.0200 3544.7900 2478.0200 3547.8100 ;
        RECT 2655.0200 3544.7900 2658.0200 3547.8100 ;
        RECT 2835.0200 3544.7900 2838.0200 3547.8100 ;
        RECT 2950.1000 3544.7900 2953.1000 3547.8100 ;
    END
# end of P/G power stripe data as pin

  END vssa1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 2917.6000 122.3800 2943.7000 125.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 122.3800 2.4000 125.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 302.3800 2943.7000 305.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 302.3800 2.4000 305.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 482.3800 2943.7000 485.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 482.3800 2.4000 485.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 662.3800 2943.7000 665.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 662.3800 2.4000 665.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 842.3800 2943.7000 845.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 842.3800 2.4000 845.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1022.3800 2943.7000 1025.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1022.3800 2.4000 1025.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1202.3800 2943.7000 1205.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1202.3800 2.4000 1205.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1382.3800 2943.7000 1385.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1382.3800 2.4000 1385.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1562.3800 2943.7000 1565.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1562.3800 2.4000 1565.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1742.3800 2943.7000 1745.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1742.3800 2.4000 1745.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1922.3800 2943.7000 1925.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1922.3800 2.4000 1925.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2102.3800 2943.7000 2105.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2102.3800 2.4000 2105.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2282.3800 2943.7000 2285.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2282.3800 2.4000 2285.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2462.3800 2943.7000 2465.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2462.3800 2.4000 2465.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2642.3800 2943.7000 2645.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2642.3800 2.4000 2645.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2822.3800 2943.7000 2825.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2822.3800 2.4000 2825.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3002.3800 2943.7000 3005.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 3002.3800 2.4000 3005.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3182.3800 2943.7000 3185.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 3182.3800 2.4000 3185.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3362.3800 2943.7000 3365.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 3362.3800 2.4000 3365.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 3535.4000 2943.7000 3538.4000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2943.7000 -18.7200 2943.7000 -15.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 117.0200 -18.7200 120.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 117.0200 3517.6000 120.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.0200 -18.7200 300.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.0200 3517.6000 300.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.0200 -18.7200 480.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.0200 3517.6000 480.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.0200 -18.7200 660.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.0200 3517.6000 660.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.0200 -18.7200 840.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.0200 3517.6000 840.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1017.0200 -18.7200 1020.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1017.0200 3517.6000 1020.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1197.0200 -18.7200 1200.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1197.0200 3517.6000 1200.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.0200 -18.7200 1380.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.0200 3517.6000 1380.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.0200 -18.7200 1560.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.0200 3517.6000 1560.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.0200 -18.7200 1740.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.0200 3517.6000 1740.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.0200 -18.7200 1920.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.0200 3517.6000 1920.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2097.0200 -18.7200 2100.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2097.0200 3517.6000 2100.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.0200 -18.7200 2280.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.0200 3517.6000 2280.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2457.0200 -18.7200 2460.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2457.0200 3517.6000 2460.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2637.0200 -18.7200 2640.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2637.0200 3517.6000 2640.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2817.0200 -18.7200 2820.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2817.0200 3517.6000 2820.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT -24.0800 3538.4000 -21.0800 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2940.7000 -18.7200 2943.7000 3538.4000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT -24.0800 -18.7200 -21.0800 3538.4000 ;
        RECT 2940.7000 -18.7200 2943.7000 3538.4000 ;
      LAYER met5 ;
        RECT -24.0800 -18.7200 2943.7000 -15.7200 ;
        RECT -24.0800 3535.4000 2943.7000 3538.4000 ;
        RECT -24.0800 -18.7300 -21.0800 -15.7100 ;
        RECT 117.0200 -18.7300 120.0200 -15.7100 ;
        RECT 297.0200 -18.7300 300.0200 -15.7100 ;
        RECT 477.0200 -18.7300 480.0200 -15.7100 ;
        RECT 1017.0200 -18.7300 1020.0200 -15.7100 ;
        RECT 657.0200 -18.7300 660.0200 -15.7100 ;
        RECT 837.0200 -18.7300 840.0200 -15.7100 ;
        RECT 1197.0200 -18.7300 1200.0200 -15.7100 ;
        RECT 1377.0200 -18.7300 1380.0200 -15.7100 ;
        RECT 1557.0200 -18.7300 1560.0200 -15.7100 ;
        RECT 1737.0200 -18.7300 1740.0200 -15.7100 ;
        RECT 1917.0200 -18.7300 1920.0200 -15.7100 ;
        RECT 2097.0200 -18.7300 2100.0200 -15.7100 ;
        RECT 2277.0200 -18.7300 2280.0200 -15.7100 ;
        RECT 2457.0200 -18.7300 2460.0200 -15.7100 ;
        RECT 2637.0200 -18.7300 2640.0200 -15.7100 ;
        RECT 2817.0200 -18.7300 2820.0200 -15.7100 ;
        RECT 2940.7000 -18.7300 2943.7000 -15.7100 ;
        RECT -24.0800 122.3700 -21.0800 125.3900 ;
        RECT -24.0800 302.3700 -21.0800 305.3900 ;
        RECT -24.0800 482.3700 -21.0800 485.3900 ;
        RECT -24.0800 662.3700 -21.0800 665.3900 ;
        RECT -24.0800 842.3700 -21.0800 845.3900 ;
        RECT -24.0800 1022.3700 -21.0800 1025.3900 ;
        RECT -24.0800 1202.3700 -21.0800 1205.3900 ;
        RECT -24.0800 1382.3700 -21.0800 1385.3900 ;
        RECT -24.0800 1562.3700 -21.0800 1565.3900 ;
        RECT -24.0800 1742.3700 -21.0800 1745.3900 ;
        RECT 2940.7000 122.3700 2943.7000 125.3900 ;
        RECT 2940.7000 302.3700 2943.7000 305.3900 ;
        RECT 2940.7000 482.3700 2943.7000 485.3900 ;
        RECT 2940.7000 662.3700 2943.7000 665.3900 ;
        RECT 2940.7000 842.3700 2943.7000 845.3900 ;
        RECT 2940.7000 1022.3700 2943.7000 1025.3900 ;
        RECT 2940.7000 1202.3700 2943.7000 1205.3900 ;
        RECT 2940.7000 1382.3700 2943.7000 1385.3900 ;
        RECT 2940.7000 1562.3700 2943.7000 1565.3900 ;
        RECT 2940.7000 1742.3700 2943.7000 1745.3900 ;
        RECT -24.0800 1922.3700 -21.0800 1925.3900 ;
        RECT -24.0800 2102.3700 -21.0800 2105.3900 ;
        RECT -24.0800 2282.3700 -21.0800 2285.3900 ;
        RECT -24.0800 2462.3700 -21.0800 2465.3900 ;
        RECT -24.0800 2642.3700 -21.0800 2645.3900 ;
        RECT -24.0800 2822.3700 -21.0800 2825.3900 ;
        RECT -24.0800 3002.3700 -21.0800 3005.3900 ;
        RECT -24.0800 3182.3700 -21.0800 3185.3900 ;
        RECT -24.0800 3362.3700 -21.0800 3365.3900 ;
        RECT 2940.7000 1922.3700 2943.7000 1925.3900 ;
        RECT 2940.7000 2102.3700 2943.7000 2105.3900 ;
        RECT 2940.7000 2282.3700 2943.7000 2285.3900 ;
        RECT 2940.7000 2462.3700 2943.7000 2465.3900 ;
        RECT 2940.7000 2642.3700 2943.7000 2645.3900 ;
        RECT 2940.7000 2822.3700 2943.7000 2825.3900 ;
        RECT 2940.7000 3002.3700 2943.7000 3005.3900 ;
        RECT 2940.7000 3182.3700 2943.7000 3185.3900 ;
        RECT 2940.7000 3362.3700 2943.7000 3365.3900 ;
        RECT -24.0800 3535.3900 -21.0800 3538.4100 ;
        RECT 117.0200 3535.3900 120.0200 3538.4100 ;
        RECT 297.0200 3535.3900 300.0200 3538.4100 ;
        RECT 477.0200 3535.3900 480.0200 3538.4100 ;
        RECT 1017.0200 3535.3900 1020.0200 3538.4100 ;
        RECT 657.0200 3535.3900 660.0200 3538.4100 ;
        RECT 837.0200 3535.3900 840.0200 3538.4100 ;
        RECT 1197.0200 3535.3900 1200.0200 3538.4100 ;
        RECT 1377.0200 3535.3900 1380.0200 3538.4100 ;
        RECT 1557.0200 3535.3900 1560.0200 3538.4100 ;
        RECT 1737.0200 3535.3900 1740.0200 3538.4100 ;
        RECT 1917.0200 3535.3900 1920.0200 3538.4100 ;
        RECT 2097.0200 3535.3900 2100.0200 3538.4100 ;
        RECT 2277.0200 3535.3900 2280.0200 3538.4100 ;
        RECT 2457.0200 3535.3900 2460.0200 3538.4100 ;
        RECT 2637.0200 3535.3900 2640.0200 3538.4100 ;
        RECT 2817.0200 3535.3900 2820.0200 3538.4100 ;
        RECT 2940.7000 3535.3900 2943.7000 3538.4100 ;
    END
# end of P/G power stripe data as pin

  END vssd2
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 2917.6000 104.1400 2934.3000 107.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 104.1400 2.4000 107.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 284.1400 2934.3000 287.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 284.1400 2.4000 287.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 464.1400 2934.3000 467.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 464.1400 2.4000 467.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 644.1400 2934.3000 647.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 644.1400 2.4000 647.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 824.1400 2934.3000 827.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 824.1400 2.4000 827.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1004.1400 2934.3000 1007.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1004.1400 2.4000 1007.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1184.1400 2934.3000 1187.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1184.1400 2.4000 1187.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1364.1400 2934.3000 1367.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1364.1400 2.4000 1367.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1544.1400 2934.3000 1547.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1544.1400 2.4000 1547.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1724.1400 2934.3000 1727.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1724.1400 2.4000 1727.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1904.1400 2934.3000 1907.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1904.1400 2.4000 1907.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2084.1400 2934.3000 2087.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2084.1400 2.4000 2087.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2264.1400 2934.3000 2267.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2264.1400 2.4000 2267.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2444.1400 2934.3000 2447.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2444.1400 2.4000 2447.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2624.1400 2934.3000 2627.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2624.1400 2.4000 2627.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2804.1400 2934.3000 2807.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2804.1400 2.4000 2807.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2984.1400 2934.3000 2987.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2984.1400 2.4000 2987.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3164.1400 2934.3000 3167.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 3164.1400 2.4000 3167.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3344.1400 2934.3000 3347.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 3344.1400 2.4000 3347.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 3526.0000 2934.3000 3529.0000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2934.3000 -9.3200 2934.3000 -6.3200 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.0200 -9.3200 102.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.0200 3517.6000 102.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 279.0200 -9.3200 282.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 279.0200 3517.6000 282.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 459.0200 -9.3200 462.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 459.0200 3517.6000 462.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 639.0200 -9.3200 642.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 639.0200 3517.6000 642.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 819.0200 -9.3200 822.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 819.0200 3517.6000 822.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 999.0200 -9.3200 1002.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 999.0200 3517.6000 1002.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1179.0200 -9.3200 1182.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1179.0200 3517.6000 1182.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1359.0200 -9.3200 1362.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1359.0200 3517.6000 1362.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1539.0200 -9.3200 1542.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1539.0200 3517.6000 1542.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.0200 -9.3200 1722.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.0200 3517.6000 1722.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1899.0200 -9.3200 1902.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1899.0200 3517.6000 1902.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2079.0200 -9.3200 2082.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2079.0200 3517.6000 2082.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2259.0200 -9.3200 2262.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2259.0200 3517.6000 2262.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2439.0200 -9.3200 2442.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2439.0200 3517.6000 2442.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2619.0200 -9.3200 2622.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2619.0200 3517.6000 2622.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2799.0200 -9.3200 2802.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2799.0200 3517.6000 2802.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT -14.6800 3529.0000 -11.6800 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.3000 -9.3200 2934.3000 3529.0000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT -14.6800 -9.3200 -11.6800 3529.0000 ;
        RECT 2931.3000 -9.3200 2934.3000 3529.0000 ;
        RECT 99.0200 0.0000 102.0200 3520.0000 ;
        RECT 279.0200 0.0000 282.0200 3520.0000 ;
        RECT 459.0200 0.0000 462.0200 3520.0000 ;
        RECT 1359.0200 323.6800 1362.0200 3520.0000 ;
        RECT 639.0200 0.0000 642.0200 3520.0000 ;
        RECT 819.0200 0.0000 822.0200 3520.0000 ;
        RECT 999.0200 0.0000 1002.0200 3520.0000 ;
        RECT 1179.0200 0.0000 1182.0200 3520.0000 ;
        RECT 1539.0200 0.0000 1542.0200 3520.0000 ;
        RECT 1719.0200 0.0000 1722.0200 3520.0000 ;
        RECT 1899.0200 0.0000 1902.0200 3520.0000 ;
        RECT 2079.0200 0.0000 2082.0200 3520.0000 ;
        RECT 2259.0200 0.0000 2262.0200 3520.0000 ;
        RECT 2439.0200 0.0000 2442.0200 3520.0000 ;
        RECT 2619.0200 0.0000 2622.0200 3520.0000 ;
        RECT 2799.0200 0.0000 2802.0200 3520.0000 ;
        RECT 1295.9200 151.2800 1299.1200 326.8800 ;
        RECT 1359.0200 0.0000 1362.0200 154.4800 ;
        RECT 1345.5350 151.2800 1348.7350 201.0000 ;
        RECT 1345.6200 151.2800 1348.8200 162.5600 ;
        RECT 1400.0200 151.2800 1403.2200 162.5600 ;
        RECT 1372.8200 151.2800 1376.0200 162.5600 ;
        RECT 1345.6200 315.6000 1348.8200 326.8800 ;
        RECT 1372.8200 315.6000 1376.0200 326.8800 ;
        RECT 1400.0200 315.6000 1403.2200 326.8800 ;
        RECT 1470.1600 151.2800 1473.3600 326.8800 ;
        RECT 1345.5350 151.2800 1348.8200 154.4800 ;
      LAYER met5 ;
        RECT -14.6800 -9.3200 2934.3000 -6.3200 ;
        RECT 0.0000 104.1400 2920.0000 107.1400 ;
        RECT 1295.9200 151.2800 1473.3600 154.4800 ;
        RECT 1295.9200 323.6800 1473.3600 326.8800 ;
        RECT 0.0000 464.1400 2920.0000 467.1400 ;
        RECT 0.0000 644.1400 2920.0000 647.1400 ;
        RECT 0.0000 824.1400 2920.0000 827.1400 ;
        RECT 0.0000 1004.1400 2920.0000 1007.1400 ;
        RECT 0.0000 1184.1400 2920.0000 1187.1400 ;
        RECT 0.0000 1364.1400 2920.0000 1367.1400 ;
        RECT 0.0000 1544.1400 2920.0000 1547.1400 ;
        RECT 0.0000 1724.1400 2920.0000 1727.1400 ;
        RECT 0.0000 284.1400 1299.1200 287.1400 ;
        RECT 1470.1600 284.1400 2920.0000 287.1400 ;
        RECT 0.0000 1904.1400 2920.0000 1907.1400 ;
        RECT 0.0000 2084.1400 2920.0000 2087.1400 ;
        RECT 0.0000 2264.1400 2920.0000 2267.1400 ;
        RECT 0.0000 2444.1400 2920.0000 2447.1400 ;
        RECT 0.0000 2624.1400 2920.0000 2627.1400 ;
        RECT 0.0000 2804.1400 2920.0000 2807.1400 ;
        RECT 0.0000 2984.1400 2920.0000 2987.1400 ;
        RECT 0.0000 3164.1400 2920.0000 3167.1400 ;
        RECT 0.0000 3344.1400 2920.0000 3347.1400 ;
        RECT -14.6800 3526.0000 2934.3000 3529.0000 ;
        RECT -14.6800 -9.3300 -11.6800 -6.3100 ;
        RECT 99.0200 -9.3300 102.0200 -6.3100 ;
        RECT 279.0200 -9.3300 282.0200 -6.3100 ;
        RECT 459.0200 -9.3300 462.0200 -6.3100 ;
        RECT 639.0200 -9.3300 642.0200 -6.3100 ;
        RECT 819.0200 -9.3300 822.0200 -6.3100 ;
        RECT 999.0200 -9.3300 1002.0200 -6.3100 ;
        RECT 1179.0200 -9.3300 1182.0200 -6.3100 ;
        RECT 1359.0200 -9.3300 1362.0200 -6.3100 ;
        RECT 1899.0200 -9.3300 1902.0200 -6.3100 ;
        RECT 1539.0200 -9.3300 1542.0200 -6.3100 ;
        RECT 1719.0200 -9.3300 1722.0200 -6.3100 ;
        RECT 2079.0200 -9.3300 2082.0200 -6.3100 ;
        RECT 2259.0200 -9.3300 2262.0200 -6.3100 ;
        RECT 2439.0200 -9.3300 2442.0200 -6.3100 ;
        RECT 2619.0200 -9.3300 2622.0200 -6.3100 ;
        RECT 2799.0200 -9.3300 2802.0200 -6.3100 ;
        RECT 2931.3000 -9.3300 2934.3000 -6.3100 ;
        RECT -14.6800 104.1300 -11.6800 107.1500 ;
        RECT -14.6800 284.1300 -11.6800 287.1500 ;
        RECT -14.6800 464.1300 -11.6800 467.1500 ;
        RECT -14.6800 644.1300 -11.6800 647.1500 ;
        RECT -14.6800 824.1300 -11.6800 827.1500 ;
        RECT -14.6800 1004.1300 -11.6800 1007.1500 ;
        RECT -14.6800 1184.1300 -11.6800 1187.1500 ;
        RECT -14.6800 1364.1300 -11.6800 1367.1500 ;
        RECT -14.6800 1544.1300 -11.6800 1547.1500 ;
        RECT -14.6800 1724.1300 -11.6800 1727.1500 ;
        RECT 2931.3000 104.1300 2934.3000 107.1500 ;
        RECT 2931.3000 284.1300 2934.3000 287.1500 ;
        RECT 2931.3000 464.1300 2934.3000 467.1500 ;
        RECT 2931.3000 644.1300 2934.3000 647.1500 ;
        RECT 2931.3000 824.1300 2934.3000 827.1500 ;
        RECT 2931.3000 1004.1300 2934.3000 1007.1500 ;
        RECT 2931.3000 1184.1300 2934.3000 1187.1500 ;
        RECT 2931.3000 1364.1300 2934.3000 1367.1500 ;
        RECT 2931.3000 1544.1300 2934.3000 1547.1500 ;
        RECT 2931.3000 1724.1300 2934.3000 1727.1500 ;
        RECT -14.6800 1904.1300 -11.6800 1907.1500 ;
        RECT -14.6800 2084.1300 -11.6800 2087.1500 ;
        RECT -14.6800 2264.1300 -11.6800 2267.1500 ;
        RECT -14.6800 2444.1300 -11.6800 2447.1500 ;
        RECT -14.6800 2624.1300 -11.6800 2627.1500 ;
        RECT -14.6800 2804.1300 -11.6800 2807.1500 ;
        RECT -14.6800 2984.1300 -11.6800 2987.1500 ;
        RECT -14.6800 3164.1300 -11.6800 3167.1500 ;
        RECT -14.6800 3344.1300 -11.6800 3347.1500 ;
        RECT 2931.3000 1904.1300 2934.3000 1907.1500 ;
        RECT 2931.3000 2084.1300 2934.3000 2087.1500 ;
        RECT 2931.3000 2264.1300 2934.3000 2267.1500 ;
        RECT 2931.3000 2444.1300 2934.3000 2447.1500 ;
        RECT 2931.3000 2624.1300 2934.3000 2627.1500 ;
        RECT 2931.3000 2804.1300 2934.3000 2807.1500 ;
        RECT 2931.3000 2984.1300 2934.3000 2987.1500 ;
        RECT 2931.3000 3164.1300 2934.3000 3167.1500 ;
        RECT 2931.3000 3344.1300 2934.3000 3347.1500 ;
        RECT -14.6800 3525.9900 -11.6800 3529.0100 ;
        RECT 99.0200 3525.9900 102.0200 3529.0100 ;
        RECT 279.0200 3525.9900 282.0200 3529.0100 ;
        RECT 459.0200 3525.9900 462.0200 3529.0100 ;
        RECT 639.0200 3525.9900 642.0200 3529.0100 ;
        RECT 819.0200 3525.9900 822.0200 3529.0100 ;
        RECT 999.0200 3525.9900 1002.0200 3529.0100 ;
        RECT 1179.0200 3525.9900 1182.0200 3529.0100 ;
        RECT 1359.0200 3525.9900 1362.0200 3529.0100 ;
        RECT 1899.0200 3525.9900 1902.0200 3529.0100 ;
        RECT 1539.0200 3525.9900 1542.0200 3529.0100 ;
        RECT 1719.0200 3525.9900 1722.0200 3529.0100 ;
        RECT 2079.0200 3525.9900 2082.0200 3529.0100 ;
        RECT 2259.0200 3525.9900 2262.0200 3529.0100 ;
        RECT 2439.0200 3525.9900 2442.0200 3529.0100 ;
        RECT 2619.0200 3525.9900 2622.0200 3529.0100 ;
        RECT 2799.0200 3525.9900 2802.0200 3529.0100 ;
        RECT 2931.3000 3525.9900 2934.3000 3529.0100 ;
    END
# end of P/G power stripe data as pin

  END vssd1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 2917.6000 68.3800 2962.5000 71.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 68.3800 2.4000 71.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 248.3800 2962.5000 251.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 248.3800 2.4000 251.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 428.3800 2962.5000 431.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 428.3800 2.4000 431.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 608.3800 2962.5000 611.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 608.3800 2.4000 611.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 788.3800 2962.5000 791.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 788.3800 2.4000 791.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 968.3800 2962.5000 971.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 968.3800 2.4000 971.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1148.3800 2962.5000 1151.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1148.3800 2.4000 1151.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1328.3800 2962.5000 1331.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1328.3800 2.4000 1331.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1508.3800 2962.5000 1511.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1508.3800 2.4000 1511.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1688.3800 2962.5000 1691.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1688.3800 2.4000 1691.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1868.3800 2962.5000 1871.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1868.3800 2.4000 1871.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2048.3800 2962.5000 2051.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2048.3800 2.4000 2051.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2228.3800 2962.5000 2231.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2228.3800 2.4000 2231.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2408.3800 2962.5000 2411.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2408.3800 2.4000 2411.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2588.3800 2962.5000 2591.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2588.3800 2.4000 2591.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2768.3800 2962.5000 2771.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2768.3800 2.4000 2771.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2948.3800 2962.5000 2951.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2948.3800 2.4000 2951.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3128.3800 2962.5000 3131.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 3128.3800 2.4000 3131.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3308.3800 2962.5000 3311.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 3308.3800 2.4000 3311.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3488.3800 2962.5000 3491.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 3488.3800 2.4000 3491.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.1800 3549.5000 2957.8000 3552.5000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2957.8000 -32.8200 2957.8000 -29.8200 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.0200 -37.5200 66.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.0200 3517.6000 66.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 243.0200 -37.5200 246.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 243.0200 3517.6000 246.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 423.0200 -37.5200 426.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 423.0200 3517.6000 426.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 603.0200 -37.5200 606.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 603.0200 3517.6000 606.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 783.0200 -37.5200 786.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 783.0200 3517.6000 786.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 963.0200 -37.5200 966.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 963.0200 3517.6000 966.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1143.0200 -37.5200 1146.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1143.0200 3517.6000 1146.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1323.0200 -37.5200 1326.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1323.0200 3517.6000 1326.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1503.0200 -37.5200 1506.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1503.0200 3517.6000 1506.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1683.0200 -37.5200 1686.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1683.0200 3517.6000 1686.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1863.0200 -37.5200 1866.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1863.0200 3517.6000 1866.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2043.0200 -37.5200 2046.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2043.0200 3517.6000 2046.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2223.0200 -37.5200 2226.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2223.0200 3517.6000 2226.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.0200 -37.5200 2406.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.0200 3517.6000 2406.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2583.0200 -37.5200 2586.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2583.0200 3517.6000 2586.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2763.0200 -37.5200 2766.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2763.0200 3517.6000 2766.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT -38.1800 3552.5000 -35.1800 3552.5000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2954.8000 -32.8200 2957.8000 3552.5000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT -38.1800 -32.8200 -35.1800 3552.5000 ;
        RECT 2954.8000 -32.8200 2957.8000 3552.5000 ;
      LAYER met5 ;
        RECT -38.1800 -32.8200 2957.8000 -29.8200 ;
        RECT -38.1800 3549.5000 2957.8000 3552.5000 ;
        RECT -38.1800 -32.8300 -35.1800 -29.8100 ;
        RECT 63.0200 -32.8300 66.0200 -29.8100 ;
        RECT 243.0200 -32.8300 246.0200 -29.8100 ;
        RECT 423.0200 -32.8300 426.0200 -29.8100 ;
        RECT 603.0200 -32.8300 606.0200 -29.8100 ;
        RECT 783.0200 -32.8300 786.0200 -29.8100 ;
        RECT 963.0200 -32.8300 966.0200 -29.8100 ;
        RECT 1143.0200 -32.8300 1146.0200 -29.8100 ;
        RECT 1323.0200 -32.8300 1326.0200 -29.8100 ;
        RECT 1503.0200 -32.8300 1506.0200 -29.8100 ;
        RECT 1683.0200 -32.8300 1686.0200 -29.8100 ;
        RECT 1863.0200 -32.8300 1866.0200 -29.8100 ;
        RECT 2043.0200 -32.8300 2046.0200 -29.8100 ;
        RECT 2223.0200 -32.8300 2226.0200 -29.8100 ;
        RECT 2403.0200 -32.8300 2406.0200 -29.8100 ;
        RECT 2763.0200 -32.8300 2766.0200 -29.8100 ;
        RECT 2583.0200 -32.8300 2586.0200 -29.8100 ;
        RECT 2954.8000 -32.8300 2957.8000 -29.8100 ;
        RECT -38.1800 68.3700 -35.1800 71.3900 ;
        RECT -38.1800 248.3700 -35.1800 251.3900 ;
        RECT -38.1800 428.3700 -35.1800 431.3900 ;
        RECT -38.1800 608.3700 -35.1800 611.3900 ;
        RECT -38.1800 788.3700 -35.1800 791.3900 ;
        RECT -38.1800 968.3700 -35.1800 971.3900 ;
        RECT -38.1800 1148.3700 -35.1800 1151.3900 ;
        RECT -38.1800 1328.3700 -35.1800 1331.3900 ;
        RECT -38.1800 1508.3700 -35.1800 1511.3900 ;
        RECT -38.1800 1688.3700 -35.1800 1691.3900 ;
        RECT 2954.8000 68.3700 2957.8000 71.3900 ;
        RECT 2954.8000 248.3700 2957.8000 251.3900 ;
        RECT 2954.8000 428.3700 2957.8000 431.3900 ;
        RECT 2954.8000 608.3700 2957.8000 611.3900 ;
        RECT 2954.8000 788.3700 2957.8000 791.3900 ;
        RECT 2954.8000 968.3700 2957.8000 971.3900 ;
        RECT 2954.8000 1148.3700 2957.8000 1151.3900 ;
        RECT 2954.8000 1328.3700 2957.8000 1331.3900 ;
        RECT 2954.8000 1508.3700 2957.8000 1511.3900 ;
        RECT 2954.8000 1688.3700 2957.8000 1691.3900 ;
        RECT -38.1800 1868.3700 -35.1800 1871.3900 ;
        RECT -38.1800 2048.3700 -35.1800 2051.3900 ;
        RECT -38.1800 2228.3700 -35.1800 2231.3900 ;
        RECT -38.1800 2408.3700 -35.1800 2411.3900 ;
        RECT -38.1800 2588.3700 -35.1800 2591.3900 ;
        RECT -38.1800 2768.3700 -35.1800 2771.3900 ;
        RECT -38.1800 2948.3700 -35.1800 2951.3900 ;
        RECT -38.1800 3128.3700 -35.1800 3131.3900 ;
        RECT -38.1800 3308.3700 -35.1800 3311.3900 ;
        RECT -38.1800 3488.3700 -35.1800 3491.3900 ;
        RECT 2954.8000 1868.3700 2957.8000 1871.3900 ;
        RECT 2954.8000 2048.3700 2957.8000 2051.3900 ;
        RECT 2954.8000 2228.3700 2957.8000 2231.3900 ;
        RECT 2954.8000 2408.3700 2957.8000 2411.3900 ;
        RECT 2954.8000 2588.3700 2957.8000 2591.3900 ;
        RECT 2954.8000 2768.3700 2957.8000 2771.3900 ;
        RECT 2954.8000 2948.3700 2957.8000 2951.3900 ;
        RECT 2954.8000 3128.3700 2957.8000 3131.3900 ;
        RECT 2954.8000 3308.3700 2957.8000 3311.3900 ;
        RECT 2954.8000 3488.3700 2957.8000 3491.3900 ;
        RECT -38.1800 3549.4900 -35.1800 3552.5100 ;
        RECT 63.0200 3549.4900 66.0200 3552.5100 ;
        RECT 243.0200 3549.4900 246.0200 3552.5100 ;
        RECT 423.0200 3549.4900 426.0200 3552.5100 ;
        RECT 603.0200 3549.4900 606.0200 3552.5100 ;
        RECT 783.0200 3549.4900 786.0200 3552.5100 ;
        RECT 963.0200 3549.4900 966.0200 3552.5100 ;
        RECT 1143.0200 3549.4900 1146.0200 3552.5100 ;
        RECT 1323.0200 3549.4900 1326.0200 3552.5100 ;
        RECT 1503.0200 3549.4900 1506.0200 3552.5100 ;
        RECT 1683.0200 3549.4900 1686.0200 3552.5100 ;
        RECT 1863.0200 3549.4900 1866.0200 3552.5100 ;
        RECT 2043.0200 3549.4900 2046.0200 3552.5100 ;
        RECT 2223.0200 3549.4900 2226.0200 3552.5100 ;
        RECT 2403.0200 3549.4900 2406.0200 3552.5100 ;
        RECT 2763.0200 3549.4900 2766.0200 3552.5100 ;
        RECT 2583.0200 3549.4900 2586.0200 3552.5100 ;
        RECT 2954.8000 3549.4900 2957.8000 3552.5100 ;
    END
# end of P/G power stripe data as pin

  END vdda2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 2917.6000 50.3800 2953.1000 53.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 50.3800 2.4000 53.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 230.3800 2953.1000 233.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 230.3800 2.4000 233.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 410.3800 2953.1000 413.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 410.3800 2.4000 413.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 590.3800 2953.1000 593.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 590.3800 2.4000 593.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 770.3800 2953.1000 773.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 770.3800 2.4000 773.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 950.3800 2953.1000 953.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 950.3800 2.4000 953.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1130.3800 2953.1000 1133.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1130.3800 2.4000 1133.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1310.3800 2953.1000 1313.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1310.3800 2.4000 1313.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1490.3800 2953.1000 1493.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1490.3800 2.4000 1493.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1670.3800 2953.1000 1673.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1670.3800 2.4000 1673.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1850.3800 2953.1000 1853.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1850.3800 2.4000 1853.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2030.3800 2953.1000 2033.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2030.3800 2.4000 2033.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2210.3800 2953.1000 2213.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2210.3800 2.4000 2213.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2390.3800 2953.1000 2393.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2390.3800 2.4000 2393.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2570.3800 2953.1000 2573.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2570.3800 2.4000 2573.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2750.3800 2953.1000 2753.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2750.3800 2.4000 2753.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2930.3800 2953.1000 2933.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2930.3800 2.4000 2933.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3110.3800 2953.1000 3113.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 3110.3800 2.4000 3113.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3290.3800 2953.1000 3293.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 3290.3800 2.4000 3293.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3470.3800 2953.1000 3473.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 3470.3800 2.4000 3473.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -28.7800 3540.1000 2948.4000 3543.1000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2948.4000 -23.4200 2948.4000 -20.4200 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.0200 -28.1200 48.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.0200 3517.6000 48.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 225.0200 -28.1200 228.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 225.0200 3517.6000 228.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.0200 -28.1200 408.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.0200 3517.6000 408.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 585.0200 -28.1200 588.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 585.0200 3517.6000 588.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 765.0200 -28.1200 768.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 765.0200 3517.6000 768.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 945.0200 -28.1200 948.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 945.0200 3517.6000 948.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1125.0200 -28.1200 1128.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1125.0200 3517.6000 1128.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1305.0200 -28.1200 1308.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1305.0200 3517.6000 1308.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1485.0200 -28.1200 1488.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1485.0200 3517.6000 1488.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1665.0200 -28.1200 1668.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1665.0200 3517.6000 1668.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1845.0200 -28.1200 1848.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1845.0200 3517.6000 1848.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2025.0200 -28.1200 2028.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2025.0200 3517.6000 2028.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2205.0200 -28.1200 2208.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2205.0200 3517.6000 2208.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2385.0200 -28.1200 2388.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2385.0200 3517.6000 2388.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2565.0200 -28.1200 2568.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2565.0200 3517.6000 2568.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2745.0200 -28.1200 2748.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2745.0200 3517.6000 2748.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT -28.7800 3543.1000 -25.7800 3543.1000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2945.4000 -23.4200 2948.4000 3543.1000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT -28.7800 -23.4200 -25.7800 3543.1000 ;
        RECT 2945.4000 -23.4200 2948.4000 3543.1000 ;
      LAYER met5 ;
        RECT -28.7800 -23.4200 2948.4000 -20.4200 ;
        RECT -28.7800 3540.1000 2948.4000 3543.1000 ;
        RECT -28.7800 -23.4300 -25.7800 -20.4100 ;
        RECT 45.0200 -23.4300 48.0200 -20.4100 ;
        RECT 225.0200 -23.4300 228.0200 -20.4100 ;
        RECT 405.0200 -23.4300 408.0200 -20.4100 ;
        RECT 585.0200 -23.4300 588.0200 -20.4100 ;
        RECT 765.0200 -23.4300 768.0200 -20.4100 ;
        RECT 945.0200 -23.4300 948.0200 -20.4100 ;
        RECT 1125.0200 -23.4300 1128.0200 -20.4100 ;
        RECT 1305.0200 -23.4300 1308.0200 -20.4100 ;
        RECT 1485.0200 -23.4300 1488.0200 -20.4100 ;
        RECT 1665.0200 -23.4300 1668.0200 -20.4100 ;
        RECT 1845.0200 -23.4300 1848.0200 -20.4100 ;
        RECT 2025.0200 -23.4300 2028.0200 -20.4100 ;
        RECT 2205.0200 -23.4300 2208.0200 -20.4100 ;
        RECT 2385.0200 -23.4300 2388.0200 -20.4100 ;
        RECT 2565.0200 -23.4300 2568.0200 -20.4100 ;
        RECT 2745.0200 -23.4300 2748.0200 -20.4100 ;
        RECT 2945.4000 -23.4300 2948.4000 -20.4100 ;
        RECT -28.7800 50.3700 -25.7800 53.3900 ;
        RECT -28.7800 230.3700 -25.7800 233.3900 ;
        RECT -28.7800 410.3700 -25.7800 413.3900 ;
        RECT -28.7800 590.3700 -25.7800 593.3900 ;
        RECT -28.7800 770.3700 -25.7800 773.3900 ;
        RECT -28.7800 950.3700 -25.7800 953.3900 ;
        RECT -28.7800 1130.3700 -25.7800 1133.3900 ;
        RECT -28.7800 1310.3700 -25.7800 1313.3900 ;
        RECT -28.7800 1490.3700 -25.7800 1493.3900 ;
        RECT -28.7800 1670.3700 -25.7800 1673.3900 ;
        RECT 2945.4000 50.3700 2948.4000 53.3900 ;
        RECT 2945.4000 230.3700 2948.4000 233.3900 ;
        RECT 2945.4000 410.3700 2948.4000 413.3900 ;
        RECT 2945.4000 590.3700 2948.4000 593.3900 ;
        RECT 2945.4000 770.3700 2948.4000 773.3900 ;
        RECT 2945.4000 950.3700 2948.4000 953.3900 ;
        RECT 2945.4000 1130.3700 2948.4000 1133.3900 ;
        RECT 2945.4000 1310.3700 2948.4000 1313.3900 ;
        RECT 2945.4000 1490.3700 2948.4000 1493.3900 ;
        RECT 2945.4000 1670.3700 2948.4000 1673.3900 ;
        RECT -28.7800 1850.3700 -25.7800 1853.3900 ;
        RECT -28.7800 2030.3700 -25.7800 2033.3900 ;
        RECT -28.7800 2210.3700 -25.7800 2213.3900 ;
        RECT -28.7800 2390.3700 -25.7800 2393.3900 ;
        RECT -28.7800 2570.3700 -25.7800 2573.3900 ;
        RECT -28.7800 2750.3700 -25.7800 2753.3900 ;
        RECT -28.7800 2930.3700 -25.7800 2933.3900 ;
        RECT -28.7800 3110.3700 -25.7800 3113.3900 ;
        RECT -28.7800 3290.3700 -25.7800 3293.3900 ;
        RECT -28.7800 3470.3700 -25.7800 3473.3900 ;
        RECT 2945.4000 1850.3700 2948.4000 1853.3900 ;
        RECT 2945.4000 2030.3700 2948.4000 2033.3900 ;
        RECT 2945.4000 2210.3700 2948.4000 2213.3900 ;
        RECT 2945.4000 2390.3700 2948.4000 2393.3900 ;
        RECT 2945.4000 2570.3700 2948.4000 2573.3900 ;
        RECT 2945.4000 2750.3700 2948.4000 2753.3900 ;
        RECT 2945.4000 2930.3700 2948.4000 2933.3900 ;
        RECT 2945.4000 3110.3700 2948.4000 3113.3900 ;
        RECT 2945.4000 3290.3700 2948.4000 3293.3900 ;
        RECT 2945.4000 3470.3700 2948.4000 3473.3900 ;
        RECT -28.7800 3540.0900 -25.7800 3543.1100 ;
        RECT 45.0200 3540.0900 48.0200 3543.1100 ;
        RECT 225.0200 3540.0900 228.0200 3543.1100 ;
        RECT 405.0200 3540.0900 408.0200 3543.1100 ;
        RECT 585.0200 3540.0900 588.0200 3543.1100 ;
        RECT 765.0200 3540.0900 768.0200 3543.1100 ;
        RECT 945.0200 3540.0900 948.0200 3543.1100 ;
        RECT 1125.0200 3540.0900 1128.0200 3543.1100 ;
        RECT 1305.0200 3540.0900 1308.0200 3543.1100 ;
        RECT 1485.0200 3540.0900 1488.0200 3543.1100 ;
        RECT 1665.0200 3540.0900 1668.0200 3543.1100 ;
        RECT 1845.0200 3540.0900 1848.0200 3543.1100 ;
        RECT 2025.0200 3540.0900 2028.0200 3543.1100 ;
        RECT 2205.0200 3540.0900 2208.0200 3543.1100 ;
        RECT 2385.0200 3540.0900 2388.0200 3543.1100 ;
        RECT 2565.0200 3540.0900 2568.0200 3543.1100 ;
        RECT 2745.0200 3540.0900 2748.0200 3543.1100 ;
        RECT 2945.4000 3540.0900 2948.4000 3543.1100 ;
    END
# end of P/G power stripe data as pin

  END vdda1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 2917.6000 32.3800 2943.7000 35.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 32.3800 2.4000 35.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 212.3800 2943.7000 215.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 212.3800 2.4000 215.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 392.3800 2943.7000 395.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 392.3800 2.4000 395.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 572.3800 2943.7000 575.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 572.3800 2.4000 575.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 752.3800 2943.7000 755.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 752.3800 2.4000 755.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 932.3800 2943.7000 935.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 932.3800 2.4000 935.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1112.3800 2943.7000 1115.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1112.3800 2.4000 1115.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1292.3800 2943.7000 1295.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1292.3800 2.4000 1295.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1472.3800 2943.7000 1475.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1472.3800 2.4000 1475.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1652.3800 2943.7000 1655.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1652.3800 2.4000 1655.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1832.3800 2943.7000 1835.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1832.3800 2.4000 1835.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2012.3800 2943.7000 2015.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2012.3800 2.4000 2015.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2192.3800 2943.7000 2195.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2192.3800 2.4000 2195.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2372.3800 2943.7000 2375.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2372.3800 2.4000 2375.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2552.3800 2943.7000 2555.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2552.3800 2.4000 2555.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2732.3800 2943.7000 2735.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2732.3800 2.4000 2735.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2912.3800 2943.7000 2915.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2912.3800 2.4000 2915.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3092.3800 2943.7000 3095.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 3092.3800 2.4000 3095.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3272.3800 2943.7000 3275.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 3272.3800 2.4000 3275.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3452.3800 2943.7000 3455.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 3452.3800 2.4000 3455.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.3800 3530.7000 2939.0000 3533.7000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2939.0000 -14.0200 2939.0000 -11.0200 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.0200 -18.7200 30.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.0200 3517.6000 30.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 207.0200 -18.7200 210.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 207.0200 3517.6000 210.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.0200 -18.7200 390.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.0200 3517.6000 390.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.0200 -18.7200 570.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.0200 3517.6000 570.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 747.0200 -18.7200 750.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 747.0200 3517.6000 750.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.0200 -18.7200 930.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.0200 3517.6000 930.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.0200 -18.7200 1110.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.0200 3517.6000 1110.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.0200 -18.7200 1290.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.0200 3517.6000 1290.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1467.0200 -18.7200 1470.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1467.0200 3517.6000 1470.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1647.0200 -18.7200 1650.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1647.0200 3517.6000 1650.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.0200 -18.7200 1830.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.0200 3517.6000 1830.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.0200 -18.7200 2010.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.0200 3517.6000 2010.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.0200 -18.7200 2190.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.0200 3517.6000 2190.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2367.0200 -18.7200 2370.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2367.0200 3517.6000 2370.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.0200 -18.7200 2550.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.0200 3517.6000 2550.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2727.0200 -18.7200 2730.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2727.0200 3517.6000 2730.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2907.0200 -18.7200 2910.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2907.0200 3517.6000 2910.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT -19.3800 3533.7000 -16.3800 3533.7000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2936.0000 -14.0200 2939.0000 3533.7000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT -19.3800 -14.0200 -16.3800 3533.7000 ;
        RECT 2936.0000 -14.0200 2939.0000 3533.7000 ;
      LAYER met5 ;
        RECT -19.3800 -14.0200 2939.0000 -11.0200 ;
        RECT -19.3800 3530.7000 2939.0000 3533.7000 ;
        RECT -19.3800 -14.0300 -16.3800 -11.0100 ;
        RECT 27.0200 -14.0300 30.0200 -11.0100 ;
        RECT 207.0200 -14.0300 210.0200 -11.0100 ;
        RECT 387.0200 -14.0300 390.0200 -11.0100 ;
        RECT 567.0200 -14.0300 570.0200 -11.0100 ;
        RECT 927.0200 -14.0300 930.0200 -11.0100 ;
        RECT 747.0200 -14.0300 750.0200 -11.0100 ;
        RECT 1287.0200 -14.0300 1290.0200 -11.0100 ;
        RECT 1107.0200 -14.0300 1110.0200 -11.0100 ;
        RECT 1827.0200 -14.0300 1830.0200 -11.0100 ;
        RECT 1647.0200 -14.0300 1650.0200 -11.0100 ;
        RECT 1467.0200 -14.0300 1470.0200 -11.0100 ;
        RECT 2187.0200 -14.0300 2190.0200 -11.0100 ;
        RECT 2007.0200 -14.0300 2010.0200 -11.0100 ;
        RECT 2727.0200 -14.0300 2730.0200 -11.0100 ;
        RECT 2547.0200 -14.0300 2550.0200 -11.0100 ;
        RECT 2367.0200 -14.0300 2370.0200 -11.0100 ;
        RECT 2936.0000 -14.0300 2939.0000 -11.0100 ;
        RECT 2907.0200 -14.0300 2910.0200 -11.0100 ;
        RECT -19.3800 32.3700 -16.3800 35.3900 ;
        RECT -19.3800 212.3700 -16.3800 215.3900 ;
        RECT -19.3800 392.3700 -16.3800 395.3900 ;
        RECT -19.3800 572.3700 -16.3800 575.3900 ;
        RECT -19.3800 752.3700 -16.3800 755.3900 ;
        RECT -19.3800 932.3700 -16.3800 935.3900 ;
        RECT -19.3800 1112.3700 -16.3800 1115.3900 ;
        RECT -19.3800 1292.3700 -16.3800 1295.3900 ;
        RECT -19.3800 1472.3700 -16.3800 1475.3900 ;
        RECT -19.3800 1652.3700 -16.3800 1655.3900 ;
        RECT 2936.0000 32.3700 2939.0000 35.3900 ;
        RECT 2936.0000 212.3700 2939.0000 215.3900 ;
        RECT 2936.0000 392.3700 2939.0000 395.3900 ;
        RECT 2936.0000 572.3700 2939.0000 575.3900 ;
        RECT 2936.0000 752.3700 2939.0000 755.3900 ;
        RECT 2936.0000 932.3700 2939.0000 935.3900 ;
        RECT 2936.0000 1112.3700 2939.0000 1115.3900 ;
        RECT 2936.0000 1292.3700 2939.0000 1295.3900 ;
        RECT 2936.0000 1472.3700 2939.0000 1475.3900 ;
        RECT 2936.0000 1652.3700 2939.0000 1655.3900 ;
        RECT -19.3800 1832.3700 -16.3800 1835.3900 ;
        RECT -19.3800 2012.3700 -16.3800 2015.3900 ;
        RECT -19.3800 2192.3700 -16.3800 2195.3900 ;
        RECT -19.3800 2372.3700 -16.3800 2375.3900 ;
        RECT -19.3800 2552.3700 -16.3800 2555.3900 ;
        RECT -19.3800 2732.3700 -16.3800 2735.3900 ;
        RECT -19.3800 2912.3700 -16.3800 2915.3900 ;
        RECT -19.3800 3092.3700 -16.3800 3095.3900 ;
        RECT -19.3800 3272.3700 -16.3800 3275.3900 ;
        RECT -19.3800 3452.3700 -16.3800 3455.3900 ;
        RECT 2936.0000 1832.3700 2939.0000 1835.3900 ;
        RECT 2936.0000 2012.3700 2939.0000 2015.3900 ;
        RECT 2936.0000 2192.3700 2939.0000 2195.3900 ;
        RECT 2936.0000 2372.3700 2939.0000 2375.3900 ;
        RECT 2936.0000 2552.3700 2939.0000 2555.3900 ;
        RECT 2936.0000 2732.3700 2939.0000 2735.3900 ;
        RECT 2936.0000 2912.3700 2939.0000 2915.3900 ;
        RECT 2936.0000 3092.3700 2939.0000 3095.3900 ;
        RECT 2936.0000 3272.3700 2939.0000 3275.3900 ;
        RECT 2936.0000 3452.3700 2939.0000 3455.3900 ;
        RECT -19.3800 3530.6900 -16.3800 3533.7100 ;
        RECT 27.0200 3530.6900 30.0200 3533.7100 ;
        RECT 207.0200 3530.6900 210.0200 3533.7100 ;
        RECT 387.0200 3530.6900 390.0200 3533.7100 ;
        RECT 567.0200 3530.6900 570.0200 3533.7100 ;
        RECT 747.0200 3530.6900 750.0200 3533.7100 ;
        RECT 927.0200 3530.6900 930.0200 3533.7100 ;
        RECT 1287.0200 3530.6900 1290.0200 3533.7100 ;
        RECT 1107.0200 3530.6900 1110.0200 3533.7100 ;
        RECT 1827.0200 3530.6900 1830.0200 3533.7100 ;
        RECT 1647.0200 3530.6900 1650.0200 3533.7100 ;
        RECT 1467.0200 3530.6900 1470.0200 3533.7100 ;
        RECT 2187.0200 3530.6900 2190.0200 3533.7100 ;
        RECT 2007.0200 3530.6900 2010.0200 3533.7100 ;
        RECT 2727.0200 3530.6900 2730.0200 3533.7100 ;
        RECT 2547.0200 3530.6900 2550.0200 3533.7100 ;
        RECT 2367.0200 3530.6900 2370.0200 3533.7100 ;
        RECT 2936.0000 3530.6900 2939.0000 3533.7100 ;
        RECT 2907.0200 3530.6900 2910.0200 3533.7100 ;
    END
# end of P/G power stripe data as pin

  END vccd2
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 2917.6000 14.1400 2934.3000 17.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 14.1400 2.4000 17.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 194.1400 2934.3000 197.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 194.1400 2.4000 197.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 374.1400 2934.3000 377.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 374.1400 2.4000 377.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 554.1400 2934.3000 557.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 554.1400 2.4000 557.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 734.1400 2934.3000 737.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 734.1400 2.4000 737.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 914.1400 2934.3000 917.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 914.1400 2.4000 917.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1094.1400 2934.3000 1097.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1094.1400 2.4000 1097.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1274.1400 2934.3000 1277.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1274.1400 2.4000 1277.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1454.1400 2934.3000 1457.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1454.1400 2.4000 1457.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1634.1400 2934.3000 1637.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1634.1400 2.4000 1637.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1814.1400 2934.3000 1817.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1814.1400 2.4000 1817.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1994.1400 2934.3000 1997.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1994.1400 2.4000 1997.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2174.1400 2934.3000 2177.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2174.1400 2.4000 2177.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2354.1400 2934.3000 2357.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2354.1400 2.4000 2357.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2534.1400 2934.3000 2537.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2534.1400 2.4000 2537.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2714.1400 2934.3000 2717.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2714.1400 2.4000 2717.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2894.1400 2934.3000 2897.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2894.1400 2.4000 2897.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3074.1400 2934.3000 3077.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 3074.1400 2.4000 3077.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3254.1400 2934.3000 3257.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 3254.1400 2.4000 3257.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3434.1400 2934.3000 3437.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 3434.1400 2.4000 3437.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.9800 3521.3000 2929.6000 3524.3000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2929.6000 -4.6200 2929.6000 -1.6200 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.0200 -9.3200 12.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.0200 3517.6000 12.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 189.0200 -9.3200 192.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 189.0200 3517.6000 192.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 369.0200 -9.3200 372.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 369.0200 3517.6000 372.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 549.0200 -9.3200 552.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 549.0200 3517.6000 552.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 729.0200 -9.3200 732.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 729.0200 3517.6000 732.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 909.0200 -9.3200 912.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 909.0200 3517.6000 912.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1089.0200 -9.3200 1092.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1089.0200 3517.6000 1092.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1269.0200 -9.3200 1272.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1269.0200 3517.6000 1272.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1449.0200 -9.3200 1452.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1449.0200 3517.6000 1452.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1629.0200 -9.3200 1632.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1629.0200 3517.6000 1632.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1809.0200 -9.3200 1812.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1809.0200 3517.6000 1812.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1989.0200 -9.3200 1992.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1989.0200 3517.6000 1992.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2169.0200 -9.3200 2172.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2169.0200 3517.6000 2172.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2349.0200 -9.3200 2352.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2349.0200 3517.6000 2352.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2529.0200 -9.3200 2532.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2529.0200 3517.6000 2532.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.0200 -9.3200 2712.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.0200 3517.6000 2712.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2889.0200 -9.3200 2892.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2889.0200 3517.6000 2892.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT -9.9800 3524.3000 -6.9800 3524.3000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2926.6000 -4.6200 2929.6000 3524.3000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT -9.9800 -4.6200 -6.9800 3524.3000 ;
        RECT 2926.6000 -4.6200 2929.6000 3524.3000 ;
        RECT 9.0200 0.0000 12.0200 3520.0000 ;
        RECT 189.0200 0.0000 192.0200 3520.0000 ;
        RECT 369.0200 0.0000 372.0200 3520.0000 ;
        RECT 549.0200 0.0000 552.0200 3520.0000 ;
        RECT 1449.0200 318.8800 1452.0200 3520.0000 ;
        RECT 729.0200 0.0000 732.0200 3520.0000 ;
        RECT 1269.0200 0.0000 1272.0200 3520.0000 ;
        RECT 1089.0200 0.0000 1092.0200 3520.0000 ;
        RECT 909.0200 0.0000 912.0200 3520.0000 ;
        RECT 1629.0200 0.0000 1632.0200 3520.0000 ;
        RECT 1809.0200 0.0000 1812.0200 3520.0000 ;
        RECT 2169.0200 0.0000 2172.0200 3520.0000 ;
        RECT 1989.0200 0.0000 1992.0200 3520.0000 ;
        RECT 2889.0200 0.0000 2892.0200 3520.0000 ;
        RECT 2709.0200 0.0000 2712.0200 3520.0000 ;
        RECT 2529.0200 0.0000 2532.0200 3520.0000 ;
        RECT 2349.0200 0.0000 2352.0200 3520.0000 ;
        RECT 1300.7200 156.0800 1303.9200 322.0800 ;
        RECT 1449.0200 0.0000 1452.0200 159.2800 ;
        RECT 1386.4200 156.0800 1389.6200 162.5600 ;
        RECT 1359.2200 156.0800 1362.4200 162.5600 ;
        RECT 1413.6200 156.0800 1416.8200 162.5600 ;
        RECT 1359.2200 315.6000 1362.4200 322.0800 ;
        RECT 1386.4200 315.6000 1389.6200 322.0800 ;
        RECT 1413.6200 315.6000 1416.8200 322.0800 ;
        RECT 1465.3600 156.0800 1468.5600 322.0800 ;
      LAYER met5 ;
        RECT -9.9800 -4.6200 2929.6000 -1.6200 ;
        RECT 0.0000 14.1400 2920.0000 17.1400 ;
        RECT 1300.7200 156.0800 1468.5600 159.2800 ;
        RECT 1300.7200 318.8800 1468.5600 322.0800 ;
        RECT 0.0000 374.1400 2920.0000 377.1400 ;
        RECT 0.0000 554.1400 2920.0000 557.1400 ;
        RECT 0.0000 734.1400 2920.0000 737.1400 ;
        RECT 0.0000 914.1400 2920.0000 917.1400 ;
        RECT 0.0000 1094.1400 2920.0000 1097.1400 ;
        RECT 0.0000 1274.1400 2920.0000 1277.1400 ;
        RECT 0.0000 1454.1400 2920.0000 1457.1400 ;
        RECT 0.0000 1634.1400 2920.0000 1637.1400 ;
        RECT 0.0000 194.1400 1303.9200 197.1400 ;
        RECT 1465.3600 194.1400 2920.0000 197.1400 ;
        RECT 0.0000 1814.1400 2920.0000 1817.1400 ;
        RECT 0.0000 1994.1400 2920.0000 1997.1400 ;
        RECT 0.0000 2174.1400 2920.0000 2177.1400 ;
        RECT 0.0000 2354.1400 2920.0000 2357.1400 ;
        RECT 0.0000 2534.1400 2920.0000 2537.1400 ;
        RECT 0.0000 2714.1400 2920.0000 2717.1400 ;
        RECT 0.0000 2894.1400 2920.0000 2897.1400 ;
        RECT 0.0000 3074.1400 2920.0000 3077.1400 ;
        RECT 0.0000 3254.1400 2920.0000 3257.1400 ;
        RECT 0.0000 3434.1400 2920.0000 3437.1400 ;
        RECT -9.9800 3521.3000 2929.6000 3524.3000 ;
        RECT 9.0200 -4.6300 12.0200 -1.6100 ;
        RECT -9.9800 -4.6300 -6.9800 -1.6100 ;
        RECT 549.0200 -4.6300 552.0200 -1.6100 ;
        RECT 369.0200 -4.6300 372.0200 -1.6100 ;
        RECT 189.0200 -4.6300 192.0200 -1.6100 ;
        RECT 909.0200 -4.6300 912.0200 -1.6100 ;
        RECT 729.0200 -4.6300 732.0200 -1.6100 ;
        RECT 1449.0200 -4.6300 1452.0200 -1.6100 ;
        RECT 1269.0200 -4.6300 1272.0200 -1.6100 ;
        RECT 1089.0200 -4.6300 1092.0200 -1.6100 ;
        RECT 1809.0200 -4.6300 1812.0200 -1.6100 ;
        RECT 1629.0200 -4.6300 1632.0200 -1.6100 ;
        RECT 2169.0200 -4.6300 2172.0200 -1.6100 ;
        RECT 1989.0200 -4.6300 1992.0200 -1.6100 ;
        RECT 2709.0200 -4.6300 2712.0200 -1.6100 ;
        RECT 2529.0200 -4.6300 2532.0200 -1.6100 ;
        RECT 2349.0200 -4.6300 2352.0200 -1.6100 ;
        RECT 2926.6000 -4.6300 2929.6000 -1.6100 ;
        RECT 2889.0200 -4.6300 2892.0200 -1.6100 ;
        RECT -9.9800 14.1300 -6.9800 17.1500 ;
        RECT -9.9800 194.1300 -6.9800 197.1500 ;
        RECT -9.9800 374.1300 -6.9800 377.1500 ;
        RECT -9.9800 554.1300 -6.9800 557.1500 ;
        RECT -9.9800 734.1300 -6.9800 737.1500 ;
        RECT -9.9800 914.1300 -6.9800 917.1500 ;
        RECT -9.9800 1094.1300 -6.9800 1097.1500 ;
        RECT -9.9800 1274.1300 -6.9800 1277.1500 ;
        RECT -9.9800 1454.1300 -6.9800 1457.1500 ;
        RECT -9.9800 1634.1300 -6.9800 1637.1500 ;
        RECT 2926.6000 14.1300 2929.6000 17.1500 ;
        RECT 2926.6000 194.1300 2929.6000 197.1500 ;
        RECT 2926.6000 374.1300 2929.6000 377.1500 ;
        RECT 2926.6000 554.1300 2929.6000 557.1500 ;
        RECT 2926.6000 734.1300 2929.6000 737.1500 ;
        RECT 2926.6000 914.1300 2929.6000 917.1500 ;
        RECT 2926.6000 1094.1300 2929.6000 1097.1500 ;
        RECT 2926.6000 1274.1300 2929.6000 1277.1500 ;
        RECT 2926.6000 1454.1300 2929.6000 1457.1500 ;
        RECT 2926.6000 1634.1300 2929.6000 1637.1500 ;
        RECT -9.9800 1814.1300 -6.9800 1817.1500 ;
        RECT -9.9800 1994.1300 -6.9800 1997.1500 ;
        RECT -9.9800 2174.1300 -6.9800 2177.1500 ;
        RECT -9.9800 2354.1300 -6.9800 2357.1500 ;
        RECT -9.9800 2534.1300 -6.9800 2537.1500 ;
        RECT -9.9800 2714.1300 -6.9800 2717.1500 ;
        RECT -9.9800 2894.1300 -6.9800 2897.1500 ;
        RECT -9.9800 3074.1300 -6.9800 3077.1500 ;
        RECT -9.9800 3254.1300 -6.9800 3257.1500 ;
        RECT -9.9800 3434.1300 -6.9800 3437.1500 ;
        RECT 2926.6000 1814.1300 2929.6000 1817.1500 ;
        RECT 2926.6000 1994.1300 2929.6000 1997.1500 ;
        RECT 2926.6000 2174.1300 2929.6000 2177.1500 ;
        RECT 2926.6000 2354.1300 2929.6000 2357.1500 ;
        RECT 2926.6000 2534.1300 2929.6000 2537.1500 ;
        RECT 2926.6000 2714.1300 2929.6000 2717.1500 ;
        RECT 2926.6000 2894.1300 2929.6000 2897.1500 ;
        RECT 2926.6000 3074.1300 2929.6000 3077.1500 ;
        RECT 2926.6000 3254.1300 2929.6000 3257.1500 ;
        RECT 2926.6000 3434.1300 2929.6000 3437.1500 ;
        RECT 9.0200 3521.2900 12.0200 3524.3100 ;
        RECT -9.9800 3521.2900 -6.9800 3524.3100 ;
        RECT 549.0200 3521.2900 552.0200 3524.3100 ;
        RECT 369.0200 3521.2900 372.0200 3524.3100 ;
        RECT 189.0200 3521.2900 192.0200 3524.3100 ;
        RECT 909.0200 3521.2900 912.0200 3524.3100 ;
        RECT 729.0200 3521.2900 732.0200 3524.3100 ;
        RECT 1449.0200 3521.2900 1452.0200 3524.3100 ;
        RECT 1269.0200 3521.2900 1272.0200 3524.3100 ;
        RECT 1089.0200 3521.2900 1092.0200 3524.3100 ;
        RECT 1809.0200 3521.2900 1812.0200 3524.3100 ;
        RECT 1629.0200 3521.2900 1632.0200 3524.3100 ;
        RECT 2169.0200 3521.2900 2172.0200 3524.3100 ;
        RECT 1989.0200 3521.2900 1992.0200 3524.3100 ;
        RECT 2709.0200 3521.2900 2712.0200 3524.3100 ;
        RECT 2529.0200 3521.2900 2532.0200 3524.3100 ;
        RECT 2349.0200 3521.2900 2352.0200 3524.3100 ;
        RECT 2926.6000 3521.2900 2929.6000 3524.3100 ;
        RECT 2889.0200 3521.2900 2892.0200 3524.3100 ;
    END
# end of P/G power stripe data as pin

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.0000 0.0000 2920.0000 3520.0000 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 2920.0000 3520.0000 ;
    LAYER met2 ;
      RECT 0.0000 0.0000 2920.0000 3520.0000 ;
    LAYER met3 ;
      RECT 0.0000 0.0000 2920.0000 3520.0000 ;
    LAYER met4 ;
      RECT 0.0000 0.0000 2920.0000 3520.0000 ;
    LAYER met5 ;
      RECT 0.0000 0.0000 2920.0000 3520.0000 ;
  END
END user_project_wrapper

END LIBRARY
