##
## LEF for PtnCells ;
## created by Innovus v17.11-s080_1 on Fri Jun 11 09:03:14 2021
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO user_project_wrapper
  CLASS BLOCK ;
  SIZE 2920.0000 BY 3520.0000 ;
  FOREIGN user_project_wrapper 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 64.708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 345.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.4503 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 147.808 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.11 LAYER met4  ;
    ANTENNAMAXAREACAR 43.0744 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 225.914 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 2.7100 -4.8000 3.2700 2.4000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.439 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.969 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 13.5102 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 66.1303 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 8.2300 -4.8000 8.7900 2.4000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.1998 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.773 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 76.8452 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 371.663 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 26.1700 -4.8000 26.7300 2.4000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.6766 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.157 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 62.546 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 308.504 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 20.1900 -4.8000 20.7500 2.4000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.289 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.875 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.504 LAYER met2  ;
    ANTENNAMAXAREACAR 48.177 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 230.367 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 32.1500 -4.8000 32.7100 2.4000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.2385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.9748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.336 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 113.658 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 582.579 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 126.4500 -4.8000 127.0100 2.4000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.2841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.1415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 6.4504 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 30.8175 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 102.9900 -4.8000 103.5500 2.4000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.2385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.9748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.336 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 107.058 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 549.579 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 79.5300 -4.8000 80.0900 2.4000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5587 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.6325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.1578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 84.8766 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 439.159 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 55.6100 -4.8000 56.1700 2.4000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.0306 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 80.045 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 79.5036 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 395.131 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 617.2700 -4.8000 617.8300 2.4000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.0404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 80.094 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 71.9295 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 357.261 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 599.3300 -4.8000 599.8900 2.4000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.381 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 76.797 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 64.4572 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 319.899 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 581.8500 -4.8000 582.4100 2.4000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.6026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 72.905 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 60.8426 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 301.826 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 563.9100 -4.8000 564.4700 2.4000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.0686 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 75.117 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 66.5606 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 329.939 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 546.4300 -4.8000 546.9900 2.4000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.6196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.872 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 56.3505 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 278.889 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 528.4900 -4.8000 529.0500 2.4000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0018 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.783 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 57.6891 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 285.055 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 511.0100 -4.8000 511.5700 2.4000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.7189 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.3155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.8898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.216 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 34.3071 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 182.042 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 493.0700 -4.8000 493.6300 2.4000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.0614 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 80.199 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 69.8592 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 346.909 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 475.5900 -4.8000 476.1500 2.4000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8382 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 83.965 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 68.9945 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 342.2 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 457.6500 -4.8000 458.2100 2.4000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.1234 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 75.509 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 86.5743 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 430.485 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 439.7100 -4.8000 440.2700 2.4000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.2666 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 71.225 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 110.179 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 548.509 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 422.2300 -4.8000 422.7900 2.4000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.6474 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.129 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 118.014 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 587.681 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 404.2900 -4.8000 404.8500 2.4000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.3618 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 71.701 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 116.022 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 577.725 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 386.8100 -4.8000 387.3700 2.4000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.133 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 66.1081 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 327.677 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 368.8700 -4.8000 369.4300 2.4000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.2716 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 76.132 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 62.8196 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 310.707 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 351.3900 -4.8000 351.9500 2.4000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.5304 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 72.534 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 60.2398 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 298.772 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 333.4500 -4.8000 334.0100 2.4000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0531 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.0945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 2.66646 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 12.5717 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 315.9700 -4.8000 316.5300 2.4000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.2934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.241 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 55.5529 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 274.901 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 298.0300 -4.8000 298.5900 2.4000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.7022 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.285 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 57.216 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 283.216 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 280.0900 -4.8000 280.6500 2.4000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.7218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.383 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 57.544 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 284.857 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 262.6100 -4.8000 263.1700 2.4000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.8178 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.863 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 48.7101 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 240.778 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 244.6700 -4.8000 245.2300 2.4000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.725 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.399 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 52.3756 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 259.105 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 227.1900 -4.8000 227.7500 2.4000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.3148 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.348 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 50.7182 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 250.818 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.2500 -4.8000 209.8100 2.4000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.2052 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.8 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 54.3158 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 268.806 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 191.7700 -4.8000 192.3300 2.4000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.4514 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.913 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 55.9311 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 276.315 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 173.8300 -4.8000 174.3900 2.4000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.358 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.446 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 53.4495 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 263.758 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 156.3500 -4.8000 156.9100 2.4000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.263 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.089 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 54.3764 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 269.018 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 138.4100 -4.8000 138.9700 2.4000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.5735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.6088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 30.384 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 29.6158 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 156.333 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 114.9500 -4.8000 115.5100 2.4000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.6296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.03 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 48.5703 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 240.424 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 91.0300 -4.8000 91.5900 2.4000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.011 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.829 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 51.1521 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 252.897 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 67.5700 -4.8000 68.1300 2.4000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.1207 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.3245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 4.21313 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 20.5152 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 43.6500 -4.8000 44.2100 2.4000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.2900 -4.8000 611.8500 2.4000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.8100 -4.8000 594.3700 2.4000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.8700 -4.8000 576.4300 2.4000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.9300 -4.8000 558.4900 2.4000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.4500 -4.8000 541.0100 2.4000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.5100 -4.8000 523.0700 2.4000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.0300 -4.8000 505.5900 2.4000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.0900 -4.8000 487.6500 2.4000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.6100 -4.8000 470.1700 2.4000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.6700 -4.8000 452.2300 2.4000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.1900 -4.8000 434.7500 2.4000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.2500 -4.8000 416.8100 2.4000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.3100 -4.8000 398.8700 2.4000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.8300 -4.8000 381.3900 2.4000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.8900 -4.8000 363.4500 2.4000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.4100 -4.8000 345.9700 2.4000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.4700 -4.8000 328.0300 2.4000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.9900 -4.8000 310.5500 2.4000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.0500 -4.8000 292.6100 2.4000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.5700 -4.8000 275.1300 2.4000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.6300 -4.8000 257.1900 2.4000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.1500 -4.8000 239.7100 2.4000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.2100 -4.8000 221.7700 2.4000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.2700 -4.8000 203.8300 2.4000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.7900 -4.8000 186.3500 2.4000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.8500 -4.8000 168.4100 2.4000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.3700 -4.8000 150.9300 2.4000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.4300 -4.8000 132.9900 2.4000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.9700 -4.8000 109.5300 2.4000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.0500 -4.8000 85.6100 2.4000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.5900 -4.8000 62.1500 2.4000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.1300 -4.8000 38.6900 2.4000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0285 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.8635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.1588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.984 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 123.756 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 639.456 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 14.2100 -4.8000 14.7700 2.4000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.9366 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.575 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 623.2500 -4.8000 623.8100 2.4000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.7134 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.341 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 605.3100 -4.8000 605.8700 2.4000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.405 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 587.8300 -4.8000 588.3900 2.4000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.271 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.247 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 569.8900 -4.8000 570.4500 2.4000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.077 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 552.4100 -4.8000 552.9700 2.4000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.3092 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.438 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 534.4700 -4.8000 535.0300 2.4000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3474 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.511 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 516.5300 -4.8000 517.0900 2.4000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.5738 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.761 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 499.0500 -4.8000 499.6100 2.4000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.2202 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 481.1100 -4.8000 481.6700 2.4000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.4586 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.185 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 463.6300 -4.8000 464.1900 2.4000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.9366 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.575 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 445.6900 -4.8000 446.2500 2.4000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.5546 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.665 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 428.2100 -4.8000 428.7700 2.4000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.5338 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.443 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 410.2700 -4.8000 410.8300 2.4000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.2206 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.995 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 392.7900 -4.8000 393.3500 2.4000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.4378 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.963 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 374.8500 -4.8000 375.4100 2.4000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.1042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.295 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 357.3700 -4.8000 357.9300 2.4000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.5538 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.661 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 339.4300 -4.8000 339.9900 2.4000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.173 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.757 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 321.4900 -4.8000 322.0500 2.4000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.7446 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.615 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 304.0100 -4.8000 304.5700 2.4000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.1738 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.761 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 286.0700 -4.8000 286.6300 2.4000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.4106 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.945 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 268.5900 -4.8000 269.1500 2.4000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.3914 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.731 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 250.6500 -4.8000 251.2100 2.4000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.1742 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.763 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 233.1700 -4.8000 233.7300 2.4000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.1978 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.645 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 215.2300 -4.8000 215.7900 2.4000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.6758 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.153 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 197.7500 -4.8000 198.3100 2.4000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.1526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.537 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 179.8100 -4.8000 180.3700 2.4000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.4862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.205 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 161.8700 -4.8000 162.4300 2.4000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.5806 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.677 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 144.3900 -4.8000 144.9500 2.4000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.1168 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.122 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 120.9300 -4.8000 121.4900 2.4000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.2902 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.225 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 97.0100 -4.8000 97.5700 2.4000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3054 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.301 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 73.5500 -4.8000 74.1100 2.4000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.343 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.489 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 49.6300 -4.8000 50.1900 2.4000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2881.3900 -4.8000 2881.9500 2.4000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2863.4500 -4.8000 2864.0100 2.4000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2845.5100 -4.8000 2846.0700 2.4000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2828.0300 -4.8000 2828.5900 2.4000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2810.0900 -4.8000 2810.6500 2.4000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2792.6100 -4.8000 2793.1700 2.4000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2774.6700 -4.8000 2775.2300 2.4000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2757.1900 -4.8000 2757.7500 2.4000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2739.2500 -4.8000 2739.8100 2.4000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2721.7700 -4.8000 2722.3300 2.4000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2703.8300 -4.8000 2704.3900 2.4000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2685.8900 -4.8000 2686.4500 2.4000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2668.4100 -4.8000 2668.9700 2.4000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2650.4700 -4.8000 2651.0300 2.4000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.9900 -4.8000 2633.5500 2.4000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2615.0500 -4.8000 2615.6100 2.4000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2597.5700 -4.8000 2598.1300 2.4000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.6300 -4.8000 2580.1900 2.4000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2562.1500 -4.8000 2562.7100 2.4000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.2100 -4.8000 2544.7700 2.4000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2526.7300 -4.8000 2527.2900 2.4000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2508.7900 -4.8000 2509.3500 2.4000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2490.8500 -4.8000 2491.4100 2.4000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.3700 -4.8000 2473.9300 2.4000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2455.4300 -4.8000 2455.9900 2.4000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.9500 -4.8000 2438.5100 2.4000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.0100 -4.8000 2420.5700 2.4000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2402.5300 -4.8000 2403.0900 2.4000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.5900 -4.8000 2385.1500 2.4000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.1100 -4.8000 2367.6700 2.4000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2349.1700 -4.8000 2349.7300 2.4000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.2300 -4.8000 2331.7900 2.4000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2313.7500 -4.8000 2314.3100 2.4000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.8100 -4.8000 2296.3700 2.4000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2278.3300 -4.8000 2278.8900 2.4000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.3900 -4.8000 2260.9500 2.4000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2242.9100 -4.8000 2243.4700 2.4000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.9700 -4.8000 2225.5300 2.4000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.4900 -4.8000 2208.0500 2.4000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.5500 -4.8000 2190.1100 2.4000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.0700 -4.8000 2172.6300 2.4000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.1300 -4.8000 2154.6900 2.4000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.1900 -4.8000 2136.7500 2.4000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.7100 -4.8000 2119.2700 2.4000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.7700 -4.8000 2101.3300 2.4000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.2900 -4.8000 2083.8500 2.4000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2065.3500 -4.8000 2065.9100 2.4000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.8700 -4.8000 2048.4300 2.4000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.9300 -4.8000 2030.4900 2.4000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.4500 -4.8000 2013.0100 2.4000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.5100 -4.8000 1995.0700 2.4000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.5700 -4.8000 1977.1300 2.4000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.0900 -4.8000 1959.6500 2.4000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.1500 -4.8000 1941.7100 2.4000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.6700 -4.8000 1924.2300 2.4000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.7300 -4.8000 1906.2900 2.4000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.2500 -4.8000 1888.8100 2.4000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.3100 -4.8000 1870.8700 2.4000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.8300 -4.8000 1853.3900 2.4000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.8900 -4.8000 1835.4500 2.4000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1817.4100 -4.8000 1817.9700 2.4000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.4700 -4.8000 1800.0300 2.4000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3438 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.493 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met2  ;
    ANTENNAMAXAREACAR 14.4052 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 67.6576 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1781.5300 -4.8000 1782.0900 2.4000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.7472 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 88.284 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.11 LAYER met2  ;
    ANTENNAMAXAREACAR 55.9434 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 278.09 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1764.0500 -4.8000 1764.6100 2.4000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.3222 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 71.267 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 60.1172 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 296.952 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1746.1100 -4.8000 1746.6700 2.4000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.0838 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 75.075 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 62.6739 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 309.735 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1728.6300 -4.8000 1729.1900 2.4000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.409 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 61.6754 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 302.418 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1710.6900 -4.8000 1711.2500 2.4000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.8162 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 78.855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 66.1586 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 325.626 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1693.2100 -4.8000 1693.7700 2.4000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.055 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.049 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 57.7952 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 286.091 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1675.2700 -4.8000 1675.8300 2.4000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.9583 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 64.6205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 3.84525 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 19.3455 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1657.7900 -4.8000 1658.3500 2.4000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.1982 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.765 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 56.1012 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 275.339 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1639.8500 -4.8000 1640.4100 2.4000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4134 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 71.841 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 59.5762 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 293.44 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1621.9100 -4.8000 1622.4700 2.4000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7298 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 61.1927 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 302.806 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1604.4300 -4.8000 1604.9900 2.4000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.0869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 75.1555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.7828 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 74.316 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 394.768 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1586.4900 -4.8000 1587.0500 2.4000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.959 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 79.569 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 74.0091 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 363.671 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1569.0100 -4.8000 1569.5700 2.4000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.1522 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 75.299 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 66.7638 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 326.806 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1551.0700 -4.8000 1551.6300 2.4000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.5654 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.601 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 52.302 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 256.616 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1533.5900 -4.8000 1534.1500 2.4000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.9192 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.37 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 57.2465 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 283.347 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1515.6500 -4.8000 1516.2100 2.4000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.7218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.383 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 56.6505 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 280.095 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1498.1700 -4.8000 1498.7300 2.4000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.4572 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.06 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 75.6954 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 373.764 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1480.2300 -4.8000 1480.7900 2.4000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.8634 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.973 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 54.223 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 267.481 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1462.7500 -4.8000 1463.3100 2.4000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.3475 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.4495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.4588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.584 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 72.1713 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 383.572 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1444.8100 -4.8000 1445.3700 2.4000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0933 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.1875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.7088 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.584 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 32.6376 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 173.244 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1426.8700 -4.8000 1427.4300 2.4000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.2938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.243 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 58.6869 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 290.277 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1409.3900 -4.8000 1409.9500 2.4000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.9999 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.7205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.1208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.448 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 21.8018 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 110.622 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1391.4500 -4.8000 1392.0100 2.4000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.7075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.3765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 232.447 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1240.18 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 5.94869 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 34.3111 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1373.9700 -4.8000 1374.5300 2.4000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.5513 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 57.5855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 3.35192 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 16.202 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1356.0300 -4.8000 1356.5900 2.4000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.5973 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.8255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 219.751 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1172.47 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 8.48606 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 45.2283 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1338.5500 -4.8000 1339.1100 2.4000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9389 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.5335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 216.439 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1154.81 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 10.9911 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 61.0747 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1320.6100 -4.8000 1321.1700 2.4000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.0491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 60.0845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 213.997 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1141.78 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.47985 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 20.224 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 34.176 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met5  ;
    ANTENNAMAXAREACAR 94.7808 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 190.723 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 1303.1300 -4.8000 1303.6900 2.4000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0086 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.817 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 46.9891 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 231.788 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1285.1900 -4.8000 1285.7500 2.4000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.6946 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.247 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 48.4598 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 239.141 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1267.2500 -4.8000 1267.8100 2.4000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.5481 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.4615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.329 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 124.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 10.6954 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 58.9455 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1249.7700 -4.8000 1250.3300 2.4000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.2805 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.2415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 196.452 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1048.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 4.85333 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 26.6222 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1231.8300 -4.8000 1232.3900 2.4000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.8834 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.191 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 39.1881 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 190.774 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1214.3500 -4.8000 1214.9100 2.4000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8242 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.895 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 41.2356 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 201.465 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1196.4100 -4.8000 1196.9700 2.4000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.9300 -4.8000 1179.4900 2.4000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.9900 -4.8000 1161.5500 2.4000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.5100 -4.8000 1144.0700 2.4000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.5700 -4.8000 1126.1300 2.4000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.6300 -4.8000 1108.1900 2.4000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.1500 -4.8000 1090.7100 2.4000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.2100 -4.8000 1072.7700 2.4000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.7300 -4.8000 1055.2900 2.4000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.7900 -4.8000 1037.3500 2.4000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.3100 -4.8000 1019.8700 2.4000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.3700 -4.8000 1001.9300 2.4000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.8900 -4.8000 984.4500 2.4000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.9500 -4.8000 966.5100 2.4000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.4700 -4.8000 949.0300 2.4000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.5300 -4.8000 931.0900 2.4000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.5900 -4.8000 913.1500 2.4000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.1100 -4.8000 895.6700 2.4000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.1700 -4.8000 877.7300 2.4000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.6900 -4.8000 860.2500 2.4000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.7500 -4.8000 842.3100 2.4000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.2700 -4.8000 824.8300 2.4000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.3300 -4.8000 806.8900 2.4000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.8500 -4.8000 789.4100 2.4000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.9100 -4.8000 771.4700 2.4000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.9700 -4.8000 753.5300 2.4000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.4900 -4.8000 736.0500 2.4000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.5500 -4.8000 718.1100 2.4000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.0700 -4.8000 700.6300 2.4000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.1300 -4.8000 682.6900 2.4000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.6500 -4.8000 665.2100 2.4000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.7100 -4.8000 647.2700 2.4000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.2300 -4.8000 629.7900 2.4000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2886.9100 -4.8000 2887.4700 2.4000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2869.4300 -4.8000 2869.9900 2.4000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2851.4900 -4.8000 2852.0500 2.4000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2834.0100 -4.8000 2834.5700 2.4000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2816.0700 -4.8000 2816.6300 2.4000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1454 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.619 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2798.5900 -4.8000 2799.1500 2.4000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2780.6500 -4.8000 2781.2100 2.4000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2763.1700 -4.8000 2763.7300 2.4000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2745.2300 -4.8000 2745.7900 2.4000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2727.2900 -4.8000 2727.8500 2.4000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.359 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2709.8100 -4.8000 2710.3700 2.4000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2691.8700 -4.8000 2692.4300 2.4000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2674.3900 -4.8000 2674.9500 2.4000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2656.4500 -4.8000 2657.0100 2.4000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2638.9700 -4.8000 2639.5300 2.4000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.941 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2621.0300 -4.8000 2621.5900 2.4000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2603.5500 -4.8000 2604.1100 2.4000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2585.6100 -4.8000 2586.1700 2.4000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2567.6700 -4.8000 2568.2300 2.4000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2550.1900 -4.8000 2550.7500 2.4000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2532.2500 -4.8000 2532.8100 2.4000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2514.7700 -4.8000 2515.3300 2.4000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3194 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.489 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2496.8300 -4.8000 2497.3900 2.4000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2479.3500 -4.8000 2479.9100 2.4000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2461.4100 -4.8000 2461.9700 2.4000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2443.9300 -4.8000 2444.4900 2.4000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2425.9900 -4.8000 2426.5500 2.4000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2408.5100 -4.8000 2409.0700 2.4000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2390.5700 -4.8000 2391.1300 2.4000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2372.6300 -4.8000 2373.1900 2.4000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2355.1500 -4.8000 2355.7100 2.4000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2337.2100 -4.8000 2337.7700 2.4000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2319.7300 -4.8000 2320.2900 2.4000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2301.7900 -4.8000 2302.3500 2.4000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2284.3100 -4.8000 2284.8700 2.4000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2266.3700 -4.8000 2266.9300 2.4000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2248.8900 -4.8000 2249.4500 2.4000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2230.9500 -4.8000 2231.5100 2.4000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2213.0100 -4.8000 2213.5700 2.4000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2195.5300 -4.8000 2196.0900 2.4000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2177.5900 -4.8000 2178.1500 2.4000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2160.1100 -4.8000 2160.6700 2.4000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2142.1700 -4.8000 2142.7300 2.4000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2124.6900 -4.8000 2125.2500 2.4000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2106.7500 -4.8000 2107.3100 2.4000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2089.2700 -4.8000 2089.8300 2.4000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2071.3300 -4.8000 2071.8900 2.4000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2053.8500 -4.8000 2054.4100 2.4000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2035.9100 -4.8000 2036.4700 2.4000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2017.9700 -4.8000 2018.5300 2.4000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2000.4900 -4.8000 2001.0500 2.4000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1982.5500 -4.8000 1983.1100 2.4000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1965.0700 -4.8000 1965.6300 2.4000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1947.1300 -4.8000 1947.6900 2.4000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1929.6500 -4.8000 1930.2100 2.4000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1911.7100 -4.8000 1912.2700 2.4000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4618 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.201 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1894.2300 -4.8000 1894.7900 2.4000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1876.2900 -4.8000 1876.8500 2.4000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1858.3500 -4.8000 1858.9100 2.4000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1840.8700 -4.8000 1841.4300 2.4000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1822.9300 -4.8000 1823.4900 2.4000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1805.4500 -4.8000 1806.0100 2.4000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4618 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.201 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1787.5100 -4.8000 1788.0700 2.4000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1770.0300 -4.8000 1770.5900 2.4000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1752.0900 -4.8000 1752.6500 2.4000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1734.6100 -4.8000 1735.1700 2.4000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1716.6700 -4.8000 1717.2300 2.4000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1699.1900 -4.8000 1699.7500 2.4000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1681.2500 -4.8000 1681.8100 2.4000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1663.3100 -4.8000 1663.8700 2.4000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1645.8300 -4.8000 1646.3900 2.4000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1627.8900 -4.8000 1628.4500 2.4000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1610.4100 -4.8000 1610.9700 2.4000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1592.4700 -4.8000 1593.0300 2.4000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1574.9900 -4.8000 1575.5500 2.4000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1557.0500 -4.8000 1557.6100 2.4000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4674 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.229 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1539.5700 -4.8000 1540.1300 2.4000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1521.6300 -4.8000 1522.1900 2.4000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1503.6900 -4.8000 1504.2500 2.4000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1486.2100 -4.8000 1486.7700 2.4000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1468.2700 -4.8000 1468.8300 2.4000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0222 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.003 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1450.7900 -4.8000 1451.3500 2.4000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1432.8500 -4.8000 1433.4100 2.4000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1415.3700 -4.8000 1415.9300 2.4000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1397.4300 -4.8000 1397.9900 2.4000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1379.9500 -4.8000 1380.5100 2.4000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1362.0100 -4.8000 1362.5700 2.4000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1344.0700 -4.8000 1344.6300 2.4000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1326.5900 -4.8000 1327.1500 2.4000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1308.6500 -4.8000 1309.2100 2.4000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1291.1700 -4.8000 1291.7300 2.4000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1273.2300 -4.8000 1273.7900 2.4000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1255.7500 -4.8000 1256.3100 2.4000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1237.8100 -4.8000 1238.3700 2.4000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1220.3300 -4.8000 1220.8900 2.4000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1202.3900 -4.8000 1202.9500 2.4000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.654 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.928 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6457 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.384 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 9.63095 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 47.6071 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.9808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 112.368 LAYER met4  ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 43.4165 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 228.554 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1184.9100 -4.8000 1185.4700 2.4000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 252.501 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1261.35 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER via2  ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.8342 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.008 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 56.403 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 217.34 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1166.9700 -4.8000 1167.5300 2.4000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.5969 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.7055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.5904 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 66.9558 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 325.384 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 161.454 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 775.855 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1149.0300 -4.8000 1149.5900 2.4000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.2997 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 76.2195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 48.2332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 225.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met3  ;
    ANTENNAMAXAREACAR 154.288 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 716.233 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.413208 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.1708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.048 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 172.691 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 815.44 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1131.5500 -4.8000 1132.1100 2.4000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6231 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.9545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 179.673 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 927.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 409.26 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2099.94 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1113.6100 -4.8000 1114.1700 2.4000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.714 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.2298 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.707 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 35.1689 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 165.952 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1096.1300 -4.8000 1096.6900 2.4000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1078.1900 -4.8000 1078.7500 2.4000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.714 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.2182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 80.983 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1060.7100 -4.8000 1061.2700 2.4000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.714 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.1176 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 95.018 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 50.1918 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 240.457 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1042.7700 -4.8000 1043.3300 2.4000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.714 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.334 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 96.208 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 49.6569 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 238.026 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1025.2900 -4.8000 1025.8500 2.4000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.714 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.6012 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 97.426 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 53.4302 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 260.703 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1007.3500 -4.8000 1007.9100 2.4000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.1738 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.761 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 989.4100 -4.8000 989.9700 2.4000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 501.573 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2492.79 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 971.9300 -4.8000 972.4900 2.4000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 498.052 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2475.13 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.9158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.688 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 953.9900 -4.8000 954.5500 2.4000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 499.122 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2480.53 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 936.5100 -4.8000 937.0700 2.4000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 506.262 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2516.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 918.5700 -4.8000 919.1300 2.4000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 502.737 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2498.61 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 901.0900 -4.8000 901.6500 2.4000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 479.107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2395.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.5124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.088 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 883.1500 -4.8000 883.7100 2.4000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 441.702 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2208.11 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.1914 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.376 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 865.6700 -4.8000 866.2300 2.4000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 44.072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 219.737 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.116 LAYER met2  ;
    ANTENNAMAXAREACAR 42.6109 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 203.599 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.443779 LAYER via2  ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.5908 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.288 LAYER met3  ;
    ANTENNAGATEAREA 1.434 LAYER met3  ;
    ANTENNAMAXAREACAR 46.5096 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 224.721 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.443779 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 847.7300 -4.8000 848.2900 2.4000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 366.742 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1833.43 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.4014 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.496 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 830.2500 -4.8000 830.8100 2.4000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 32.8256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 163.45 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.434 LAYER met2  ;
    ANTENNAMAXAREACAR 26.0108 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 120.684 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 812.3100 -4.8000 812.8700 2.4000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.1511 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3567 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.168 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 29.9462 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 147.392 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.815487 LAYER via3  ;
    ANTENNADIFFAREA 0.429 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.9158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.688 LAYER met4  ;
    ANTENNAGATEAREA 1.434 LAYER met4  ;
    ANTENNAMAXAREACAR 37.5583 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 188.318 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.815487 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 794.3700 -4.8000 794.9300 2.4000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.4761 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.2195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 63.6987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 340.192 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 159.118 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 834.349 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.498027 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 776.8900 -4.8000 777.4500 2.4000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.6502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 92.799 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 49.0697 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 239.98 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 758.9500 -4.8000 759.5100 2.4000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.2041 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 85.4245 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 58.7553 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 287.552 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.358176 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 59.6445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 293.354 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 741.4700 -4.8000 742.0300 2.4000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6863 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.0445 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 80.4103 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 388.536 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.41 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.32 LAYER met3  ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 123.347 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 621.234 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via3  ;
    ANTENNADIFFAREA 0.43675 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.5467 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 110.048 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 169.623 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 869.09 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 723.5300 -4.8000 724.0900 2.4000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.2508 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 85.694 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 44.9651 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 214.346 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 706.0500 -4.8000 706.6100 2.4000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8303 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 83.6465 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 41.0259 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 195.095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.498027 LAYER via2  ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.0868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.6 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 52.4827 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 257.258 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.498027 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 688.1100 -4.8000 688.6700 2.4000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.7362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 83.111 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 63.7441 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 307.362 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 670.6300 -4.8000 671.1900 2.4000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.5904 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 54.5783 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 272.269 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met2  ;
    ANTENNAMAXAREACAR 130.78 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 647.118 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.498027 LAYER via2  ;
    ANTENNADIFFAREA 1.5904 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.8604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.944 LAYER met3  ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 186.772 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 872.217 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.498027 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 652.6900 -4.8000 653.2500 2.4000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.9826 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 109.473 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 45.0586 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 208.12 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.109 LAYER met3  ;
    ANTENNAMAXAREACAR 97.1188 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 459.534 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.761465 LAYER via3  ;
    ANTENNADIFFAREA 1.5904 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.0858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.928 LAYER met4  ;
    ANTENNAGATEAREA 1.109 LAYER met4  ;
    ANTENNAMAXAREACAR 105.312 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 503.653 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.761465 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 634.7500 -4.8000 635.3100 2.4000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2892.8900 -4.8000 2893.4500 2.4000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2875.4100 -4.8000 2875.9700 2.4000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2857.4700 -4.8000 2858.0300 2.4000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2839.9900 -4.8000 2840.5500 2.4000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2822.0500 -4.8000 2822.6100 2.4000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2804.1100 -4.8000 2804.6700 2.4000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2786.6300 -4.8000 2787.1900 2.4000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2768.6900 -4.8000 2769.2500 2.4000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2751.2100 -4.8000 2751.7700 2.4000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2733.2700 -4.8000 2733.8300 2.4000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2715.7900 -4.8000 2716.3500 2.4000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2697.8500 -4.8000 2698.4100 2.4000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2680.3700 -4.8000 2680.9300 2.4000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2662.4300 -4.8000 2662.9900 2.4000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2644.9500 -4.8000 2645.5100 2.4000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2627.0100 -4.8000 2627.5700 2.4000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.0700 -4.8000 2609.6300 2.4000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2591.5900 -4.8000 2592.1500 2.4000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2573.6500 -4.8000 2574.2100 2.4000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2556.1700 -4.8000 2556.7300 2.4000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.2300 -4.8000 2538.7900 2.4000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2520.7500 -4.8000 2521.3100 2.4000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2502.8100 -4.8000 2503.3700 2.4000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.3300 -4.8000 2485.8900 2.4000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2467.3900 -4.8000 2467.9500 2.4000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2449.4500 -4.8000 2450.0100 2.4000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.9700 -4.8000 2432.5300 2.4000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2414.0300 -4.8000 2414.5900 2.4000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.5500 -4.8000 2397.1100 2.4000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.6100 -4.8000 2379.1700 2.4000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.1300 -4.8000 2361.6900 2.4000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2343.1900 -4.8000 2343.7500 2.4000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2325.7100 -4.8000 2326.2700 2.4000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2307.7700 -4.8000 2308.3300 2.4000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.2900 -4.8000 2290.8500 2.4000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2272.3500 -4.8000 2272.9100 2.4000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2254.4100 -4.8000 2254.9700 2.4000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2236.9300 -4.8000 2237.4900 2.4000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.9900 -4.8000 2219.5500 2.4000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.5100 -4.8000 2202.0700 2.4000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.5700 -4.8000 2184.1300 2.4000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2166.0900 -4.8000 2166.6500 2.4000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.1500 -4.8000 2148.7100 2.4000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.6700 -4.8000 2131.2300 2.4000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.7300 -4.8000 2113.2900 2.4000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.7900 -4.8000 2095.3500 2.4000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.3100 -4.8000 2077.8700 2.4000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.3700 -4.8000 2059.9300 2.4000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.8900 -4.8000 2042.4500 2.4000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2023.9500 -4.8000 2024.5100 2.4000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.4700 -4.8000 2007.0300 2.4000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.5300 -4.8000 1989.0900 2.4000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.0500 -4.8000 1971.6100 2.4000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.1100 -4.8000 1953.6700 2.4000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.6300 -4.8000 1936.1900 2.4000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.6900 -4.8000 1918.2500 2.4000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.7500 -4.8000 1900.3100 2.4000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.2700 -4.8000 1882.8300 2.4000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.3300 -4.8000 1864.8900 2.4000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.8500 -4.8000 1847.4100 2.4000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.9100 -4.8000 1829.4700 2.4000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1811.4300 -4.8000 1811.9900 2.4000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.861 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.16 LAYER met2  ;
    ANTENNAMAXAREACAR 7.24751 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 33.8793 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.103838 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1793.4900 -4.8000 1794.0500 2.4000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9162 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.355 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.33 LAYER met2  ;
    ANTENNAMAXAREACAR 4.72286 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.7831 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0386466 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1776.0100 -4.8000 1776.5700 2.4000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.5318 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.433 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 51.4788 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 255.158 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1758.0700 -4.8000 1758.6300 2.4000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.9414 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.363 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 58.6646 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 288.394 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1740.1300 -4.8000 1740.6900 2.4000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.327 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.409 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 55.8954 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 274.131 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1722.6500 -4.8000 1723.2100 2.4000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.675 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.149 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 50.0012 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 244.661 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1704.7100 -4.8000 1705.2700 2.4000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.6082 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.697 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 57.3305 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 283.667 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1687.2300 -4.8000 1687.7900 2.4000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.0558 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 60.053 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 50.7325 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 247.424 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1669.2900 -4.8000 1669.8500 2.4000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.904 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.294 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 41.8368 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 203.218 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1651.8100 -4.8000 1652.3700 2.4000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.8038 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.793 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 49.4808 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 242.059 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1633.8700 -4.8000 1634.4300 2.4000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.3754 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.651 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 47.9834 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 233.679 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1616.3900 -4.8000 1616.9500 2.4000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.3968 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.758 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 45.3281 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 224.131 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1598.4500 -4.8000 1599.0100 2.4000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.2462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.005 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 50.5265 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 250.123 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1580.9700 -4.8000 1581.5300 2.4000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.151 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 60.529 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 50.9224 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 252.103 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1563.0300 -4.8000 1563.5900 2.4000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.6044 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.796 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 40.8545 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 198.927 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1545.0900 -4.8000 1545.6500 2.4000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.7399 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.4205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 4.42505 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 20.0566 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1527.6100 -4.8000 1528.1700 2.4000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.3112 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.212 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 42.7083 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 210.556 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1509.6700 -4.8000 1510.2300 2.4000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.7746 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.529 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 45.101 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 222.519 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1492.1900 -4.8000 1492.7500 2.4000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.9832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.69 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 34.5644 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 167.477 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1474.2500 -4.8000 1474.8100 2.4000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.1207 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.3245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 3.38465 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 17.3414 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1456.7700 -4.8000 1457.3300 2.4000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.959 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 50.3406 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 246.358 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1438.8300 -4.8000 1439.3900 2.4000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.8868 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.208 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 45.0339 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 222.661 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1421.3500 -4.8000 1421.9100 2.4000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.2791 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.2245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 3.12566 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 16.2101 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1403.4100 -4.8000 1403.9700 2.4000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7219 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.4385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 5.01495 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 23.3212 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1385.4700 -4.8000 1386.0300 2.4000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.1042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.295 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 43.1341 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 210.325 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1367.9900 -4.8000 1368.5500 2.4000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.581 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.679 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 36.9531 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 178.527 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1350.0500 -4.8000 1350.6100 2.4000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.133 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 35.0747 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 173.137 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1332.5700 -4.8000 1333.1300 2.4000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8186 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.867 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 53.6214 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 262.762 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1314.6300 -4.8000 1315.1900 2.4000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.1979 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.8185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 4.30505 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 21.9879 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1297.1500 -4.8000 1297.7100 2.4000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9134 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.341 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 52.6218 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 256.871 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1279.2100 -4.8000 1279.7700 2.4000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.8182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.865 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 57.7281 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 283.295 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1261.7300 -4.8000 1262.2900 2.4000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6331 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.0045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 195.463 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1042.94 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 8.91434 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 50.1253 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1243.7900 -4.8000 1244.3500 2.4000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0487 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.9645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 145.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met4  ;
    ANTENNAMAXAREACAR 8.77252 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 49.2364 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1225.8500 -4.8000 1226.4100 2.4000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.0098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.823 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 33.2081 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 163.804 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1208.3700 -4.8000 1208.9300 2.4000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.4300 -4.8000 1190.9900 2.4000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.9500 -4.8000 1173.5100 2.4000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.0100 -4.8000 1155.5700 2.4000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.5300 -4.8000 1138.0900 2.4000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.5900 -4.8000 1120.1500 2.4000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.1100 -4.8000 1102.6700 2.4000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.1700 -4.8000 1084.7300 2.4000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.6900 -4.8000 1067.2500 2.4000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.7500 -4.8000 1049.3100 2.4000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.8100 -4.8000 1031.3700 2.4000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.3300 -4.8000 1013.8900 2.4000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.3900 -4.8000 995.9500 2.4000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.9100 -4.8000 978.4700 2.4000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.9700 -4.8000 960.5300 2.4000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.4900 -4.8000 943.0500 2.4000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.5500 -4.8000 925.1100 2.4000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.0700 -4.8000 907.6300 2.4000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.1300 -4.8000 889.6900 2.4000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.1900 -4.8000 871.7500 2.4000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.7100 -4.8000 854.2700 2.4000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.7700 -4.8000 836.3300 2.4000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.2900 -4.8000 818.8500 2.4000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.3500 -4.8000 800.9100 2.4000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.8700 -4.8000 783.4300 2.4000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.9300 -4.8000 765.4900 2.4000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.4500 -4.8000 748.0100 2.4000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.5100 -4.8000 730.0700 2.4000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.0300 -4.8000 712.5900 2.4000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.0900 -4.8000 694.6500 2.4000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.1500 -4.8000 676.7100 2.4000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.6700 -4.8000 659.2300 2.4000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.7300 -4.8000 641.2900 2.4000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 161.5800 2.4000 162.7800 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 357.4200 2.4000 358.6200 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 552.5800 2.4000 553.7800 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 813.7000 2.4000 814.9000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1074.1400 2.4000 1075.3400 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1335.2600 2.4000 1336.4600 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1595.7000 2.4000 1596.9000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1856.1400 2.4000 1857.3400 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2117.2600 2.4000 2118.4600 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2377.7000 2.4000 2378.9000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2638.8200 2.4000 2640.0200 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2899.2600 2.4000 2900.4600 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 3159.7000 2.4000 3160.9000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 3420.8200 2.4000 3422.0200 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.3500 3517.6000 202.9100 3524.8000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.1100 3517.6000 527.6700 3524.8000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.4100 3517.6000 851.9700 3524.8000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.7100 3517.6000 1176.2700 3524.8000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.4700 3517.6000 1501.0300 3524.8000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.7700 3517.6000 1825.3300 3524.8000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.0700 3517.6000 2149.6300 3524.8000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.8300 3517.6000 2474.3900 3524.8000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.1300 3517.6000 2798.6900 3524.8000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 3352.8200 2924.8000 3354.0200 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 3086.9400 2924.8000 3088.1400 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2821.0600 2924.8000 2822.2600 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2555.8600 2924.8000 2557.0600 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2289.9800 2924.8000 2291.1800 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2024.1000 2924.8000 2025.3000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1758.9000 2924.8000 1760.1000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1493.0200 2924.8000 1494.2200 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1227.1400 2924.8000 1228.3400 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1027.9000 2924.8000 1029.1000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 828.6600 2924.8000 829.8600 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 629.4200 2924.8000 630.6200 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 430.1800 2924.8000 431.3800 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 230.9400 2924.8000 232.1400 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 32.3800 2924.8000 33.5800 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.00495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.024 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 96.3000 2.4000 97.5000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 292.1400 2.4000 293.3400 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.8244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 487.3000 2.4000 488.5000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.8244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 748.4200 2.4000 749.6200 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.8244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1008.8600 2.4000 1010.0600 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1269.9800 2.4000 1271.1800 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.6724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met3  ;
    ANTENNAMAXAREACAR 417.712 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2089.03 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.346263 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.9808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 112.368 LAYER met4  ;
    ANTENNAGATEAREA 0.621 LAYER met4  ;
    ANTENNAMAXAREACAR 451.497 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2269.98 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.346263 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1530.4200 2.4000 1531.6200 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.1942 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.568 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 31.9689 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 172.45 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1791.5400 2.4000 1792.7400 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.5904 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 58.3158 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 311.944 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 131.342 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 702.577 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2051.9800 2.4000 2053.1800 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 39.5932 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 211.616 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met3  ;
    ANTENNAMAXAREACAR 124.507 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 665.459 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.125786 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.1708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.048 LAYER met4  ;
    ANTENNAGATEAREA 0.444 LAYER met4  ;
    ANTENNAMAXAREACAR 142.91 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 764.666 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.125786 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2312.4200 2.4000 2313.6200 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 171.033 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 913.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 385.209 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2057.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2573.5400 2.4000 2574.7400 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0752 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.0114 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.056 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2833.9800 2.4000 2835.1800 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0752 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.5324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.168 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 3095.1000 2.4000 3096.3000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.6504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.464 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 3355.5400 2.4000 3356.7400 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0752 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 404.753 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2023.54 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 121.3900 3517.6000 121.9500 3524.8000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0752 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 414.977 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2074.78 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 445.6900 3517.6000 446.2500 3524.8000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0752 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 414.151 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2070.65 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 770.4500 3517.6000 771.0100 3524.8000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0752 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 415.796 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2078.75 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1094.7500 3517.6000 1095.3100 3524.8000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 501.546 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2492.56 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1419.0500 3517.6000 1419.6100 3524.8000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 498.025 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2474.9 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.9158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.688 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1743.8100 3517.6000 1744.3700 3524.8000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 499.095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2480.3 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2068.1100 3517.6000 2068.6700 3524.8000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 506.236 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2515.89 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2392.4100 3517.6000 2392.9700 3524.8000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 502.711 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2498.38 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2717.1700 3517.6000 2717.7300 3524.8000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.8724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.648 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 3418.7800 2924.8000 3419.9800 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5514 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.936 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 3153.5800 2924.8000 3154.7800 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.07095 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2887.7000 2924.8000 2888.9000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.7614 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.056 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2621.8200 2924.8000 2623.0200 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.6564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.496 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2356.6200 2924.8000 2357.8200 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2090.7400 2924.8000 2091.9400 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0752 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.3164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1824.8600 2924.8000 1826.0600 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0752 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.6644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1559.6600 2924.8000 1560.8600 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0752 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.3164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1293.7800 2924.8000 1294.9800 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0752 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1094.5400 2924.8000 1095.7400 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0752 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.2204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 895.3000 2924.8000 896.5000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0752 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.3164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 696.0600 2924.8000 697.2600 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0752 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.0804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.424 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 496.8200 2924.8000 498.0200 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.5904 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.2204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.444 LAYER met3  ;
    ANTENNAMAXAREACAR 36.5324 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 194.829 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 297.5800 2924.8000 298.7800 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 36.4186 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 194.68 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.109 LAYER met3  ;
    ANTENNAMAXAREACAR 32.8391 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 175.546 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.0360685 LAYER via3  ;
    ANTENNADIFFAREA 1.5904 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.0858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.928 LAYER met4  ;
    ANTENNAGATEAREA 1.109 LAYER met4  ;
    ANTENNAMAXAREACAR 41.0319 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 219.665 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0360685 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 98.3400 2924.8000 99.5400 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.088 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 31.7000 2.4000 32.9000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.0004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 605.735 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3231.02 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 226.8600 2.4000 228.0600 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 605.735 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3231.02 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 422.7000 2.4000 423.9000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 605.735 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3231.02 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 683.1400 2.4000 684.3400 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 605.735 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3231.02 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 943.5800 2.4000 944.7800 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0152 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 605.735 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3231.02 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1204.7000 2.4000 1205.9000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0038 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 605.735 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3231.02 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1465.1400 2.4000 1466.3400 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 605.735 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3231.02 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1726.2600 2.4000 1727.4600 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0076 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 605.735 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3231.02 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1986.7000 2.4000 1987.9000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3886 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 605.735 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3231.02 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2247.1400 2.4000 2248.3400 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.12 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met3  ;
    ANTENNAMAXAREACAR 321.095 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1608.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.132727 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 156.584 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 835.584 LAYER met4  ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 479.261 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2452.1 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.132727 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2508.2600 2.4000 2509.4600 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.4422 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met3  ;
    ANTENNAMAXAREACAR 30.7497 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 98.5293 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2768.7000 2.4000 2769.9000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.98 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 156.584 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 835.584 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 158.165 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 844.024 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 3029.8200 2.4000 3031.0200 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 145.928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 648.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 279.117 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1489.09 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT -4.8000 3290.2600 2.4000 3291.4600 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 73.1365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 350.675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.521 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 156.584 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 835.584 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 158.165 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 844.024 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 40.4300 3517.6000 40.9900 3524.8000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 273.26 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1320.86 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 154.439 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 660.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 279.117 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1489.09 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 364.7300 3517.6000 365.2900 3524.8000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 73.1071 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 350.43 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.521 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 156.584 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 835.584 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met4  ;
    ANTENNAMAXAREACAR 158.165 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 844.024 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 689.0300 3517.6000 689.5900 3524.8000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 273.26 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1320.86 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 154.439 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 660.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 279.117 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1489.09 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1013.7900 3517.6000 1014.3500 3524.8000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 125.451 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 597.132 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.6854 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 697.945 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3723.3 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1338.0900 3517.6000 1338.6500 3524.8000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 273.26 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1320.86 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 154.439 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 660.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 279.117 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1489.09 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1662.3900 3517.6000 1662.9500 3524.8000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 125.451 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 597.132 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.6854 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 697.945 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3723.3 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1987.1500 3517.6000 1987.7100 3524.8000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 273.23 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1320.61 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 154.439 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 660.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 279.117 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1489.09 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2311.4500 3517.6000 2312.0100 3524.8000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 125.412 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 596.838 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.6854 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 697.945 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3723.3 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2635.7500 3517.6000 2636.3100 3524.8000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 145.922 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 648.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 279.117 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1489.09 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 3485.4200 2924.8000 3486.6200 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.17545 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 697.945 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3723.3 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 3219.5400 2924.8000 3220.7400 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 145.922 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 648.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 279.117 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1489.09 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2954.3400 2924.8000 2955.5400 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0454 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 697.945 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3723.3 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2688.4600 2924.8000 2689.6600 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 145.922 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 648.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 279.117 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1489.09 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2422.5800 2924.8000 2423.7800 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2866 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 697.945 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3723.3 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2157.3800 2924.8000 2158.5800 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 145.799 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 647 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 279.117 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1489.09 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1891.5000 2924.8000 1892.7000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9076 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 697.945 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3723.3 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1625.6200 2924.8000 1626.8200 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0494 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 279.117 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1489.09 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1360.4200 2924.8000 1361.6200 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9076 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 697.945 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3723.3 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1161.1800 2924.8000 1162.3800 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.6988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 279.117 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1489.09 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 961.9400 2924.8000 963.1400 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2236 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 697.945 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3723.3 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 762.7000 2924.8000 763.9000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.4662 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.672 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met3  ;
    ANTENNAMAXAREACAR 57.9503 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 232.356 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0923232 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 563.4600 2924.8000 564.6600 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.673 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 697.945 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3723.3 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 364.2200 2924.8000 365.4200 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.3432 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.536 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met3  ;
    ANTENNAMAXAREACAR 30.6497 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 97.5111 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 164.9800 2924.8000 166.1800 ;
    END
  END io_oeb[0]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 617.8600 2.4000 619.0600 ;
    END
  END analog_io[28]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 878.9800 2.4000 880.1800 ;
    END
  END analog_io[27]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1139.4200 2.4000 1140.6200 ;
    END
  END analog_io[26]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1399.8600 2.4000 1401.0600 ;
    END
  END analog_io[25]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1660.9800 2.4000 1662.1800 ;
    END
  END analog_io[24]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 1921.4200 2.4000 1922.6200 ;
    END
  END analog_io[23]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2182.5400 2.4000 2183.7400 ;
    END
  END analog_io[22]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2442.9800 2.4000 2444.1800 ;
    END
  END analog_io[21]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2703.4200 2.4000 2704.6200 ;
    END
  END analog_io[20]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 2964.5400 2.4000 2965.7400 ;
    END
  END analog_io[19]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 3224.9800 2.4000 3226.1800 ;
    END
  END analog_io[18]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.8000 3486.1000 2.4000 3487.3000 ;
    END
  END analog_io[17]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.7700 3517.6000 284.3300 3524.8000 ;
    END
  END analog_io[16]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.0700 3517.6000 608.6300 3524.8000 ;
    END
  END analog_io[15]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.3700 3517.6000 932.9300 3524.8000 ;
    END
  END analog_io[14]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.1300 3517.6000 1257.6900 3524.8000 ;
    END
  END analog_io[13]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.4300 3517.6000 1581.9900 3524.8000 ;
    END
  END analog_io[12]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.7300 3517.6000 1906.2900 3524.8000 ;
    END
  END analog_io[11]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.4900 3517.6000 2231.0500 3524.8000 ;
    END
  END analog_io[10]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.7900 3517.6000 2555.3500 3524.8000 ;
    END
  END analog_io[9]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.0900 3517.6000 2879.6500 3524.8000 ;
    END
  END analog_io[8]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 3286.1800 2924.8000 3287.3800 ;
    END
  END analog_io[7]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 3020.3000 2924.8000 3021.5000 ;
    END
  END analog_io[6]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2755.1000 2924.8000 2756.3000 ;
    END
  END analog_io[5]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2489.2200 2924.8000 2490.4200 ;
    END
  END analog_io[4]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 2223.3400 2924.8000 2224.5400 ;
    END
  END analog_io[3]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1958.1400 2924.8000 1959.3400 ;
    END
  END analog_io[2]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1692.2600 2924.8000 1693.4600 ;
    END
  END analog_io[1]
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.6000 1426.3800 2924.8000 1427.5800 ;
    END
  END analog_io[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.8700 -4.8000 2899.4300 2.4000 ;
    END
  END user_clock2
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2234 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.009 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2916.8100 -4.8000 2917.3700 2.4000 ;
    END
  END user_irq[2]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4618 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.201 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2910.8300 -4.8000 2911.3900 2.4000 ;
    END
  END user_irq[1]
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.43675 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7002 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.393 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2904.8500 -4.8000 2905.4100 2.4000 ;
    END
  END user_irq[0]
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 2917.6000 158.3800 2962.5000 161.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 158.3800 2.4000 161.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 338.3800 2962.5000 341.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 338.3800 2.4000 341.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 518.3800 2962.5000 521.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 518.3800 2.4000 521.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 698.3800 2962.5000 701.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 698.3800 2.4000 701.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 878.3800 2962.5000 881.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 878.3800 2.4000 881.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1058.3800 2962.5000 1061.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1058.3800 2.4000 1061.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1238.3800 2962.5000 1241.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1238.3800 2.4000 1241.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1418.3800 2962.5000 1421.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1418.3800 2.4000 1421.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1598.3800 2962.5000 1601.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1598.3800 2.4000 1601.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1778.3800 2962.5000 1781.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1778.3800 2.4000 1781.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1958.3800 2962.5000 1961.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1958.3800 2.4000 1961.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2138.3800 2962.5000 2141.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2138.3800 2.4000 2141.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2318.3800 2962.5000 2321.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2318.3800 2.4000 2321.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2498.3800 2962.5000 2501.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2498.3800 2.4000 2501.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2678.3800 2962.5000 2681.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2678.3800 2.4000 2681.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2858.3800 2962.5000 2861.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2858.3800 2.4000 2861.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3038.3800 2962.5000 3041.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 3038.3800 2.4000 3041.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3218.3800 2962.5000 3221.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 3218.3800 2.4000 3221.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3398.3800 2962.5000 3401.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 3398.3800 2.4000 3401.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 3554.2000 2962.5000 3557.2000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2962.5000 -37.5200 2962.5000 -34.5200 ;
    END
    PORT
      LAYER met4 ;
        RECT 153.0200 -37.5200 156.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 153.0200 3517.6000 156.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 333.0200 -37.5200 336.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 333.0200 3517.6000 336.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 513.0200 -37.5200 516.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 513.0200 3517.6000 516.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.0200 -37.5200 696.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 693.0200 3517.6000 696.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 873.0200 -37.5200 876.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 873.0200 3517.6000 876.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.0200 -37.5200 1056.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.0200 3517.6000 1056.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1233.0200 -37.5200 1236.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1233.0200 3517.6000 1236.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1413.0200 -37.5200 1416.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1413.0200 3517.6000 1416.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1593.0200 -37.5200 1596.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1593.0200 3517.6000 1596.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1773.0200 -37.5200 1776.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1773.0200 3517.6000 1776.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1953.0200 -37.5200 1956.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1953.0200 3517.6000 1956.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2133.0200 -37.5200 2136.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2133.0200 3517.6000 2136.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2313.0200 -37.5200 2316.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2313.0200 3517.6000 2316.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2493.0200 -37.5200 2496.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2493.0200 3517.6000 2496.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2673.0200 -37.5200 2676.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2673.0200 3517.6000 2676.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2853.0200 -37.5200 2856.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2853.0200 3517.6000 2856.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT -42.8800 3557.2000 -39.8800 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2959.5000 -37.5200 2962.5000 3557.2000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT 2959.5000 -37.5200 2962.5000 3557.2000 ;
        RECT -42.8800 -37.5200 -39.8800 3557.2000 ;
      LAYER met5 ;
        RECT -42.8800 -37.5200 2962.5000 -34.5200 ;
        RECT -42.8800 3554.2000 2962.5000 3557.2000 ;
        RECT -42.8800 -37.5300 -39.8800 -34.5100 ;
        RECT 513.0200 -37.5300 516.0200 -34.5100 ;
        RECT 333.0200 -37.5300 336.0200 -34.5100 ;
        RECT 153.0200 -37.5300 156.0200 -34.5100 ;
        RECT 873.0200 -37.5300 876.0200 -34.5100 ;
        RECT 693.0200 -37.5300 696.0200 -34.5100 ;
        RECT 1413.0200 -37.5300 1416.0200 -34.5100 ;
        RECT 1233.0200 -37.5300 1236.0200 -34.5100 ;
        RECT 1053.0200 -37.5300 1056.0200 -34.5100 ;
        RECT 1773.0200 -37.5300 1776.0200 -34.5100 ;
        RECT 1593.0200 -37.5300 1596.0200 -34.5100 ;
        RECT 2313.0200 -37.5300 2316.0200 -34.5100 ;
        RECT 2133.0200 -37.5300 2136.0200 -34.5100 ;
        RECT 1953.0200 -37.5300 1956.0200 -34.5100 ;
        RECT 2673.0200 -37.5300 2676.0200 -34.5100 ;
        RECT 2493.0200 -37.5300 2496.0200 -34.5100 ;
        RECT 2959.5000 -37.5300 2962.5000 -34.5100 ;
        RECT 2853.0200 -37.5300 2856.0200 -34.5100 ;
        RECT -42.8800 878.3700 -39.8800 881.3900 ;
        RECT -42.8800 158.3700 -39.8800 161.3900 ;
        RECT -42.8800 338.3700 -39.8800 341.3900 ;
        RECT -42.8800 518.3700 -39.8800 521.3900 ;
        RECT -42.8800 698.3700 -39.8800 701.3900 ;
        RECT -42.8800 1058.3700 -39.8800 1061.3900 ;
        RECT -42.8800 1238.3700 -39.8800 1241.3900 ;
        RECT -42.8800 1418.3700 -39.8800 1421.3900 ;
        RECT -42.8800 1598.3700 -39.8800 1601.3900 ;
        RECT 2959.5000 878.3700 2962.5000 881.3900 ;
        RECT 2959.5000 158.3700 2962.5000 161.3900 ;
        RECT 2959.5000 338.3700 2962.5000 341.3900 ;
        RECT 2959.5000 518.3700 2962.5000 521.3900 ;
        RECT 2959.5000 698.3700 2962.5000 701.3900 ;
        RECT 2959.5000 1058.3700 2962.5000 1061.3900 ;
        RECT 2959.5000 1238.3700 2962.5000 1241.3900 ;
        RECT 2959.5000 1418.3700 2962.5000 1421.3900 ;
        RECT 2959.5000 1598.3700 2962.5000 1601.3900 ;
        RECT -42.8800 1778.3700 -39.8800 1781.3900 ;
        RECT -42.8800 1958.3700 -39.8800 1961.3900 ;
        RECT -42.8800 2138.3700 -39.8800 2141.3900 ;
        RECT -42.8800 2318.3700 -39.8800 2321.3900 ;
        RECT -42.8800 2498.3700 -39.8800 2501.3900 ;
        RECT -42.8800 2858.3700 -39.8800 2861.3900 ;
        RECT -42.8800 2678.3700 -39.8800 2681.3900 ;
        RECT -42.8800 3038.3700 -39.8800 3041.3900 ;
        RECT -42.8800 3218.3700 -39.8800 3221.3900 ;
        RECT -42.8800 3398.3700 -39.8800 3401.3900 ;
        RECT 2959.5000 1778.3700 2962.5000 1781.3900 ;
        RECT 2959.5000 1958.3700 2962.5000 1961.3900 ;
        RECT 2959.5000 2138.3700 2962.5000 2141.3900 ;
        RECT 2959.5000 2318.3700 2962.5000 2321.3900 ;
        RECT 2959.5000 2498.3700 2962.5000 2501.3900 ;
        RECT 2959.5000 2858.3700 2962.5000 2861.3900 ;
        RECT 2959.5000 2678.3700 2962.5000 2681.3900 ;
        RECT 2959.5000 3038.3700 2962.5000 3041.3900 ;
        RECT 2959.5000 3218.3700 2962.5000 3221.3900 ;
        RECT 2959.5000 3398.3700 2962.5000 3401.3900 ;
        RECT -42.8800 3554.1900 -39.8800 3557.2100 ;
        RECT 513.0200 3554.1900 516.0200 3557.2100 ;
        RECT 333.0200 3554.1900 336.0200 3557.2100 ;
        RECT 153.0200 3554.1900 156.0200 3557.2100 ;
        RECT 873.0200 3554.1900 876.0200 3557.2100 ;
        RECT 693.0200 3554.1900 696.0200 3557.2100 ;
        RECT 1413.0200 3554.1900 1416.0200 3557.2100 ;
        RECT 1233.0200 3554.1900 1236.0200 3557.2100 ;
        RECT 1053.0200 3554.1900 1056.0200 3557.2100 ;
        RECT 1773.0200 3554.1900 1776.0200 3557.2100 ;
        RECT 1593.0200 3554.1900 1596.0200 3557.2100 ;
        RECT 2313.0200 3554.1900 2316.0200 3557.2100 ;
        RECT 2133.0200 3554.1900 2136.0200 3557.2100 ;
        RECT 1953.0200 3554.1900 1956.0200 3557.2100 ;
        RECT 2673.0200 3554.1900 2676.0200 3557.2100 ;
        RECT 2493.0200 3554.1900 2496.0200 3557.2100 ;
        RECT 2959.5000 3554.1900 2962.5000 3557.2100 ;
        RECT 2853.0200 3554.1900 2856.0200 3557.2100 ;
    END
# end of P/G power stripe data as pin

  END vssa2
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 2917.6000 140.3800 2953.1000 143.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 140.3800 2.4000 143.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 320.3800 2953.1000 323.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 320.3800 2.4000 323.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 500.3800 2953.1000 503.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 500.3800 2.4000 503.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 680.3800 2953.1000 683.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 680.3800 2.4000 683.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 860.3800 2953.1000 863.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 860.3800 2.4000 863.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1040.3800 2953.1000 1043.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1040.3800 2.4000 1043.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1220.3800 2953.1000 1223.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1220.3800 2.4000 1223.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1400.3800 2953.1000 1403.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1400.3800 2.4000 1403.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1580.3800 2953.1000 1583.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1580.3800 2.4000 1583.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1760.3800 2953.1000 1763.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1760.3800 2.4000 1763.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1940.3800 2953.1000 1943.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1940.3800 2.4000 1943.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2120.3800 2953.1000 2123.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2120.3800 2.4000 2123.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2300.3800 2953.1000 2303.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2300.3800 2.4000 2303.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2480.3800 2953.1000 2483.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2480.3800 2.4000 2483.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2660.3800 2953.1000 2663.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2660.3800 2.4000 2663.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2840.3800 2953.1000 2843.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2840.3800 2.4000 2843.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3020.3800 2953.1000 3023.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 3020.3800 2.4000 3023.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3200.3800 2953.1000 3203.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 3200.3800 2.4000 3203.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3380.3800 2953.1000 3383.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 3380.3800 2.4000 3383.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 3544.8000 2953.1000 3547.8000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2953.1000 -28.1200 2953.1000 -25.1200 ;
    END
    PORT
      LAYER met4 ;
        RECT 135.0200 -28.1200 138.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 135.0200 3517.6000 138.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 315.0200 -28.1200 318.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 315.0200 3517.6000 318.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 495.0200 -28.1200 498.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 495.0200 3517.6000 498.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.0200 -28.1200 678.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.0200 3517.6000 678.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 855.0200 -28.1200 858.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 855.0200 3517.6000 858.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1035.0200 -28.1200 1038.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1035.0200 3517.6000 1038.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1215.0200 -28.1200 1218.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1215.0200 3517.6000 1218.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1395.0200 -28.1200 1398.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1395.0200 3517.6000 1398.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1575.0200 -28.1200 1578.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1575.0200 3517.6000 1578.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1755.0200 -28.1200 1758.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1755.0200 3517.6000 1758.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1935.0200 -28.1200 1938.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1935.0200 3517.6000 1938.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2115.0200 -28.1200 2118.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2115.0200 3517.6000 2118.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2295.0200 -28.1200 2298.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2295.0200 3517.6000 2298.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2475.0200 -28.1200 2478.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2475.0200 3517.6000 2478.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2655.0200 -28.1200 2658.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2655.0200 3517.6000 2658.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2835.0200 -28.1200 2838.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2835.0200 3517.6000 2838.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT -33.4800 3547.8000 -30.4800 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2950.1000 -28.1200 2953.1000 3547.8000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT 2950.1000 -28.1200 2953.1000 3547.8000 ;
        RECT -33.4800 -28.1200 -30.4800 3547.8000 ;
      LAYER met5 ;
        RECT -33.4800 -28.1200 2953.1000 -25.1200 ;
        RECT -33.4800 3544.8000 2953.1000 3547.8000 ;
        RECT 135.0200 -28.1300 138.0200 -25.1100 ;
        RECT -33.4800 -28.1300 -30.4800 -25.1100 ;
        RECT 495.0200 -28.1300 498.0200 -25.1100 ;
        RECT 315.0200 -28.1300 318.0200 -25.1100 ;
        RECT 855.0200 -28.1300 858.0200 -25.1100 ;
        RECT 675.0200 -28.1300 678.0200 -25.1100 ;
        RECT 1215.0200 -28.1300 1218.0200 -25.1100 ;
        RECT 1395.0200 -28.1300 1398.0200 -25.1100 ;
        RECT 1035.0200 -28.1300 1038.0200 -25.1100 ;
        RECT 1755.0200 -28.1300 1758.0200 -25.1100 ;
        RECT 1575.0200 -28.1300 1578.0200 -25.1100 ;
        RECT 2115.0200 -28.1300 2118.0200 -25.1100 ;
        RECT 2295.0200 -28.1300 2298.0200 -25.1100 ;
        RECT 1935.0200 -28.1300 1938.0200 -25.1100 ;
        RECT 2655.0200 -28.1300 2658.0200 -25.1100 ;
        RECT 2475.0200 -28.1300 2478.0200 -25.1100 ;
        RECT 2950.1000 -28.1300 2953.1000 -25.1100 ;
        RECT 2835.0200 -28.1300 2838.0200 -25.1100 ;
        RECT -33.4800 140.3700 -30.4800 143.3900 ;
        RECT -33.4800 320.3700 -30.4800 323.3900 ;
        RECT -33.4800 500.3700 -30.4800 503.3900 ;
        RECT -33.4800 680.3700 -30.4800 683.3900 ;
        RECT -33.4800 860.3700 -30.4800 863.3900 ;
        RECT -33.4800 1040.3700 -30.4800 1043.3900 ;
        RECT -33.4800 1220.3700 -30.4800 1223.3900 ;
        RECT -33.4800 1400.3700 -30.4800 1403.3900 ;
        RECT -33.4800 1580.3700 -30.4800 1583.3900 ;
        RECT 2950.1000 140.3700 2953.1000 143.3900 ;
        RECT 2950.1000 320.3700 2953.1000 323.3900 ;
        RECT 2950.1000 500.3700 2953.1000 503.3900 ;
        RECT 2950.1000 680.3700 2953.1000 683.3900 ;
        RECT 2950.1000 860.3700 2953.1000 863.3900 ;
        RECT 2950.1000 1040.3700 2953.1000 1043.3900 ;
        RECT 2950.1000 1220.3700 2953.1000 1223.3900 ;
        RECT 2950.1000 1400.3700 2953.1000 1403.3900 ;
        RECT 2950.1000 1580.3700 2953.1000 1583.3900 ;
        RECT -33.4800 1760.3700 -30.4800 1763.3900 ;
        RECT -33.4800 1940.3700 -30.4800 1943.3900 ;
        RECT -33.4800 2120.3700 -30.4800 2123.3900 ;
        RECT -33.4800 2300.3700 -30.4800 2303.3900 ;
        RECT -33.4800 2480.3700 -30.4800 2483.3900 ;
        RECT -33.4800 2660.3700 -30.4800 2663.3900 ;
        RECT -33.4800 2840.3700 -30.4800 2843.3900 ;
        RECT -33.4800 3020.3700 -30.4800 3023.3900 ;
        RECT -33.4800 3200.3700 -30.4800 3203.3900 ;
        RECT -33.4800 3380.3700 -30.4800 3383.3900 ;
        RECT 2950.1000 1760.3700 2953.1000 1763.3900 ;
        RECT 2950.1000 1940.3700 2953.1000 1943.3900 ;
        RECT 2950.1000 2120.3700 2953.1000 2123.3900 ;
        RECT 2950.1000 2300.3700 2953.1000 2303.3900 ;
        RECT 2950.1000 2480.3700 2953.1000 2483.3900 ;
        RECT 2950.1000 2660.3700 2953.1000 2663.3900 ;
        RECT 2950.1000 2840.3700 2953.1000 2843.3900 ;
        RECT 2950.1000 3020.3700 2953.1000 3023.3900 ;
        RECT 2950.1000 3200.3700 2953.1000 3203.3900 ;
        RECT 2950.1000 3380.3700 2953.1000 3383.3900 ;
        RECT 135.0200 3544.7900 138.0200 3547.8100 ;
        RECT -33.4800 3544.7900 -30.4800 3547.8100 ;
        RECT 495.0200 3544.7900 498.0200 3547.8100 ;
        RECT 315.0200 3544.7900 318.0200 3547.8100 ;
        RECT 855.0200 3544.7900 858.0200 3547.8100 ;
        RECT 675.0200 3544.7900 678.0200 3547.8100 ;
        RECT 1215.0200 3544.7900 1218.0200 3547.8100 ;
        RECT 1395.0200 3544.7900 1398.0200 3547.8100 ;
        RECT 1035.0200 3544.7900 1038.0200 3547.8100 ;
        RECT 1755.0200 3544.7900 1758.0200 3547.8100 ;
        RECT 1575.0200 3544.7900 1578.0200 3547.8100 ;
        RECT 2115.0200 3544.7900 2118.0200 3547.8100 ;
        RECT 2295.0200 3544.7900 2298.0200 3547.8100 ;
        RECT 1935.0200 3544.7900 1938.0200 3547.8100 ;
        RECT 2655.0200 3544.7900 2658.0200 3547.8100 ;
        RECT 2475.0200 3544.7900 2478.0200 3547.8100 ;
        RECT 2950.1000 3544.7900 2953.1000 3547.8100 ;
        RECT 2835.0200 3544.7900 2838.0200 3547.8100 ;
    END
# end of P/G power stripe data as pin

  END vssa1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 2917.6000 122.3800 2943.7000 125.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 122.3800 2.4000 125.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 302.3800 2943.7000 305.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 302.3800 2.4000 305.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 482.3800 2943.7000 485.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 482.3800 2.4000 485.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 662.3800 2943.7000 665.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 662.3800 2.4000 665.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 842.3800 2943.7000 845.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 842.3800 2.4000 845.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1022.3800 2943.7000 1025.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1022.3800 2.4000 1025.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1202.3800 2943.7000 1205.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1202.3800 2.4000 1205.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1382.3800 2943.7000 1385.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1382.3800 2.4000 1385.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1562.3800 2943.7000 1565.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1562.3800 2.4000 1565.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1742.3800 2943.7000 1745.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1742.3800 2.4000 1745.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1922.3800 2943.7000 1925.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1922.3800 2.4000 1925.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2102.3800 2943.7000 2105.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2102.3800 2.4000 2105.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2282.3800 2943.7000 2285.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2282.3800 2.4000 2285.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2462.3800 2943.7000 2465.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2462.3800 2.4000 2465.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2642.3800 2943.7000 2645.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2642.3800 2.4000 2645.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2822.3800 2943.7000 2825.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2822.3800 2.4000 2825.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3002.3800 2943.7000 3005.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 3002.3800 2.4000 3005.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3182.3800 2943.7000 3185.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 3182.3800 2.4000 3185.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3362.3800 2943.7000 3365.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 3362.3800 2.4000 3365.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 3535.4000 2943.7000 3538.4000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2943.7000 -18.7200 2943.7000 -15.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 117.0200 -18.7200 120.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 117.0200 3517.6000 120.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.0200 -18.7200 300.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.0200 3517.6000 300.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.0200 -18.7200 480.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.0200 3517.6000 480.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.0200 -18.7200 660.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.0200 3517.6000 660.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.0200 -18.7200 840.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.0200 3517.6000 840.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1017.0200 -18.7200 1020.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1017.0200 3517.6000 1020.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1197.0200 -18.7200 1200.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1197.0200 3517.6000 1200.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.0200 -18.7200 1380.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.0200 3517.6000 1380.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.0200 -18.7200 1560.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.0200 3517.6000 1560.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.0200 -18.7200 1740.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.0200 3517.6000 1740.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.0200 -18.7200 1920.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.0200 3517.6000 1920.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2097.0200 -18.7200 2100.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2097.0200 3517.6000 2100.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.0200 -18.7200 2280.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.0200 3517.6000 2280.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2457.0200 -18.7200 2460.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2457.0200 3517.6000 2460.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2637.0200 -18.7200 2640.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2637.0200 3517.6000 2640.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2817.0200 -18.7200 2820.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2817.0200 3517.6000 2820.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT -24.0800 3538.4000 -21.0800 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2940.7000 -18.7200 2943.7000 3538.4000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT 2940.7000 -18.7200 2943.7000 3538.4000 ;
        RECT -24.0800 -18.7200 -21.0800 3538.4000 ;
      LAYER met5 ;
        RECT -24.0800 -18.7200 2943.7000 -15.7200 ;
        RECT -24.0800 3535.4000 2943.7000 3538.4000 ;
        RECT 117.0200 -18.7300 120.0200 -15.7100 ;
        RECT -24.0800 -18.7300 -21.0800 -15.7100 ;
        RECT 477.0200 -18.7300 480.0200 -15.7100 ;
        RECT 297.0200 -18.7300 300.0200 -15.7100 ;
        RECT 1017.0200 -18.7300 1020.0200 -15.7100 ;
        RECT 837.0200 -18.7300 840.0200 -15.7100 ;
        RECT 657.0200 -18.7300 660.0200 -15.7100 ;
        RECT 1377.0200 -18.7300 1380.0200 -15.7100 ;
        RECT 1197.0200 -18.7300 1200.0200 -15.7100 ;
        RECT 1737.0200 -18.7300 1740.0200 -15.7100 ;
        RECT 1557.0200 -18.7300 1560.0200 -15.7100 ;
        RECT 2277.0200 -18.7300 2280.0200 -15.7100 ;
        RECT 2097.0200 -18.7300 2100.0200 -15.7100 ;
        RECT 1917.0200 -18.7300 1920.0200 -15.7100 ;
        RECT 2637.0200 -18.7300 2640.0200 -15.7100 ;
        RECT 2457.0200 -18.7300 2460.0200 -15.7100 ;
        RECT 2940.7000 -18.7300 2943.7000 -15.7100 ;
        RECT 2817.0200 -18.7300 2820.0200 -15.7100 ;
        RECT -24.0800 122.3700 -21.0800 125.3900 ;
        RECT -24.0800 302.3700 -21.0800 305.3900 ;
        RECT -24.0800 482.3700 -21.0800 485.3900 ;
        RECT -24.0800 662.3700 -21.0800 665.3900 ;
        RECT -24.0800 842.3700 -21.0800 845.3900 ;
        RECT -24.0800 1022.3700 -21.0800 1025.3900 ;
        RECT -24.0800 1202.3700 -21.0800 1205.3900 ;
        RECT -24.0800 1382.3700 -21.0800 1385.3900 ;
        RECT -24.0800 1562.3700 -21.0800 1565.3900 ;
        RECT -24.0800 1742.3700 -21.0800 1745.3900 ;
        RECT 2940.7000 122.3700 2943.7000 125.3900 ;
        RECT 2940.7000 302.3700 2943.7000 305.3900 ;
        RECT 2940.7000 482.3700 2943.7000 485.3900 ;
        RECT 2940.7000 662.3700 2943.7000 665.3900 ;
        RECT 2940.7000 842.3700 2943.7000 845.3900 ;
        RECT 2940.7000 1022.3700 2943.7000 1025.3900 ;
        RECT 2940.7000 1202.3700 2943.7000 1205.3900 ;
        RECT 2940.7000 1382.3700 2943.7000 1385.3900 ;
        RECT 2940.7000 1562.3700 2943.7000 1565.3900 ;
        RECT 2940.7000 1742.3700 2943.7000 1745.3900 ;
        RECT -24.0800 1922.3700 -21.0800 1925.3900 ;
        RECT -24.0800 2102.3700 -21.0800 2105.3900 ;
        RECT -24.0800 2282.3700 -21.0800 2285.3900 ;
        RECT -24.0800 2462.3700 -21.0800 2465.3900 ;
        RECT -24.0800 2642.3700 -21.0800 2645.3900 ;
        RECT -24.0800 2822.3700 -21.0800 2825.3900 ;
        RECT -24.0800 3002.3700 -21.0800 3005.3900 ;
        RECT -24.0800 3182.3700 -21.0800 3185.3900 ;
        RECT -24.0800 3362.3700 -21.0800 3365.3900 ;
        RECT 2940.7000 1922.3700 2943.7000 1925.3900 ;
        RECT 2940.7000 2102.3700 2943.7000 2105.3900 ;
        RECT 2940.7000 2282.3700 2943.7000 2285.3900 ;
        RECT 2940.7000 2462.3700 2943.7000 2465.3900 ;
        RECT 2940.7000 2642.3700 2943.7000 2645.3900 ;
        RECT 2940.7000 2822.3700 2943.7000 2825.3900 ;
        RECT 2940.7000 3002.3700 2943.7000 3005.3900 ;
        RECT 2940.7000 3182.3700 2943.7000 3185.3900 ;
        RECT 2940.7000 3362.3700 2943.7000 3365.3900 ;
        RECT 117.0200 3535.3900 120.0200 3538.4100 ;
        RECT -24.0800 3535.3900 -21.0800 3538.4100 ;
        RECT 477.0200 3535.3900 480.0200 3538.4100 ;
        RECT 297.0200 3535.3900 300.0200 3538.4100 ;
        RECT 1017.0200 3535.3900 1020.0200 3538.4100 ;
        RECT 837.0200 3535.3900 840.0200 3538.4100 ;
        RECT 657.0200 3535.3900 660.0200 3538.4100 ;
        RECT 1377.0200 3535.3900 1380.0200 3538.4100 ;
        RECT 1197.0200 3535.3900 1200.0200 3538.4100 ;
        RECT 1737.0200 3535.3900 1740.0200 3538.4100 ;
        RECT 1557.0200 3535.3900 1560.0200 3538.4100 ;
        RECT 2277.0200 3535.3900 2280.0200 3538.4100 ;
        RECT 2097.0200 3535.3900 2100.0200 3538.4100 ;
        RECT 1917.0200 3535.3900 1920.0200 3538.4100 ;
        RECT 2637.0200 3535.3900 2640.0200 3538.4100 ;
        RECT 2457.0200 3535.3900 2460.0200 3538.4100 ;
        RECT 2940.7000 3535.3900 2943.7000 3538.4100 ;
        RECT 2817.0200 3535.3900 2820.0200 3538.4100 ;
    END
# end of P/G power stripe data as pin

  END vssd2
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 2917.6000 104.1400 2934.3000 107.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 104.1400 2.4000 107.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 284.1400 2934.3000 287.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 284.1400 2.4000 287.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 464.1400 2934.3000 467.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 464.1400 2.4000 467.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 644.1400 2934.3000 647.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 644.1400 2.4000 647.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 824.1400 2934.3000 827.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 824.1400 2.4000 827.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1004.1400 2934.3000 1007.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1004.1400 2.4000 1007.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1184.1400 2934.3000 1187.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1184.1400 2.4000 1187.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1364.1400 2934.3000 1367.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1364.1400 2.4000 1367.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1544.1400 2934.3000 1547.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1544.1400 2.4000 1547.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1724.1400 2934.3000 1727.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1724.1400 2.4000 1727.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1904.1400 2934.3000 1907.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1904.1400 2.4000 1907.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2084.1400 2934.3000 2087.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2084.1400 2.4000 2087.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2264.1400 2934.3000 2267.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2264.1400 2.4000 2267.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2444.1400 2934.3000 2447.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2444.1400 2.4000 2447.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2624.1400 2934.3000 2627.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2624.1400 2.4000 2627.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2804.1400 2934.3000 2807.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2804.1400 2.4000 2807.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2984.1400 2934.3000 2987.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2984.1400 2.4000 2987.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3164.1400 2934.3000 3167.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 3164.1400 2.4000 3167.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3344.1400 2934.3000 3347.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 3344.1400 2.4000 3347.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 3526.0000 2934.3000 3529.0000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2934.3000 -9.3200 2934.3000 -6.3200 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.0200 -9.3200 102.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.0200 3517.6000 102.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 279.0200 -9.3200 282.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 279.0200 3517.6000 282.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 459.0200 -9.3200 462.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 459.0200 3517.6000 462.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 639.0200 -9.3200 642.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 639.0200 3517.6000 642.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 819.0200 -9.3200 822.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 819.0200 3517.6000 822.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 999.0200 -9.3200 1002.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 999.0200 3517.6000 1002.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1179.0200 -9.3200 1182.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1179.0200 3517.6000 1182.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1359.0200 -9.3200 1362.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1359.0200 3517.6000 1362.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1539.0200 -9.3200 1542.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1539.0200 3517.6000 1542.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.0200 -9.3200 1722.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1719.0200 3517.6000 1722.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1899.0200 -9.3200 1902.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1899.0200 3517.6000 1902.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2079.0200 -9.3200 2082.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2079.0200 3517.6000 2082.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2259.0200 -9.3200 2262.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2259.0200 3517.6000 2262.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2439.0200 -9.3200 2442.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2439.0200 3517.6000 2442.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2619.0200 -9.3200 2622.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2619.0200 3517.6000 2622.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2799.0200 -9.3200 2802.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2799.0200 3517.6000 2802.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT -14.6800 3529.0000 -11.6800 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.3000 -9.3200 2934.3000 3529.0000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT 2931.3000 -9.3200 2934.3000 3529.0000 ;
        RECT -14.6800 -9.3200 -11.6800 3529.0000 ;
        RECT 459.0200 0.0000 462.0200 3520.0000 ;
        RECT 279.0200 0.0000 282.0200 3520.0000 ;
        RECT 99.0200 0.0000 102.0200 3520.0000 ;
        RECT 1359.0200 0.0000 1362.0200 3520.0000 ;
        RECT 1179.0200 0.0000 1182.0200 3520.0000 ;
        RECT 999.0200 0.0000 1002.0200 3520.0000 ;
        RECT 819.0200 0.0000 822.0200 3520.0000 ;
        RECT 639.0200 0.0000 642.0200 3520.0000 ;
        RECT 2259.0200 0.0000 2262.0200 3520.0000 ;
        RECT 2079.0200 0.0000 2082.0200 3520.0000 ;
        RECT 1899.0200 0.0000 1902.0200 3520.0000 ;
        RECT 1719.0200 0.0000 1722.0200 3520.0000 ;
        RECT 1539.0200 0.0000 1542.0200 3520.0000 ;
        RECT 2799.0200 0.0000 2802.0200 3520.0000 ;
        RECT 2619.0200 0.0000 2622.0200 3520.0000 ;
        RECT 2439.0200 0.0000 2442.0200 3520.0000 ;
      LAYER met5 ;
        RECT -14.6800 -9.3200 2934.3000 -6.3200 ;
        RECT 0.0000 104.1400 2920.0000 107.1400 ;
        RECT 0.0000 284.1400 2920.0000 287.1400 ;
        RECT 0.0000 464.1400 2920.0000 467.1400 ;
        RECT 0.0000 644.1400 2920.0000 647.1400 ;
        RECT 0.0000 824.1400 2920.0000 827.1400 ;
        RECT 0.0000 1004.1400 2920.0000 1007.1400 ;
        RECT 0.0000 1184.1400 2920.0000 1187.1400 ;
        RECT 0.0000 1364.1400 2920.0000 1367.1400 ;
        RECT 0.0000 1544.1400 2920.0000 1547.1400 ;
        RECT 0.0000 1724.1400 2920.0000 1727.1400 ;
        RECT 0.0000 1904.1400 2920.0000 1907.1400 ;
        RECT 0.0000 2084.1400 2920.0000 2087.1400 ;
        RECT 0.0000 2264.1400 2920.0000 2267.1400 ;
        RECT 0.0000 2444.1400 2920.0000 2447.1400 ;
        RECT 0.0000 2624.1400 2920.0000 2627.1400 ;
        RECT 0.0000 2804.1400 2920.0000 2807.1400 ;
        RECT 0.0000 2984.1400 2920.0000 2987.1400 ;
        RECT 0.0000 3164.1400 2920.0000 3167.1400 ;
        RECT 0.0000 3344.1400 2920.0000 3347.1400 ;
        RECT -14.6800 3526.0000 2934.3000 3529.0000 ;
        RECT 99.0200 -9.3300 102.0200 -6.3100 ;
        RECT -14.6800 -9.3300 -11.6800 -6.3100 ;
        RECT 459.0200 -9.3300 462.0200 -6.3100 ;
        RECT 279.0200 -9.3300 282.0200 -6.3100 ;
        RECT 999.0200 -9.3300 1002.0200 -6.3100 ;
        RECT 819.0200 -9.3300 822.0200 -6.3100 ;
        RECT 639.0200 -9.3300 642.0200 -6.3100 ;
        RECT 1359.0200 -9.3300 1362.0200 -6.3100 ;
        RECT 1179.0200 -9.3300 1182.0200 -6.3100 ;
        RECT 1899.0200 -9.3300 1902.0200 -6.3100 ;
        RECT 1719.0200 -9.3300 1722.0200 -6.3100 ;
        RECT 1539.0200 -9.3300 1542.0200 -6.3100 ;
        RECT 2259.0200 -9.3300 2262.0200 -6.3100 ;
        RECT 2079.0200 -9.3300 2082.0200 -6.3100 ;
        RECT 2619.0200 -9.3300 2622.0200 -6.3100 ;
        RECT 2439.0200 -9.3300 2442.0200 -6.3100 ;
        RECT 2931.3000 -9.3300 2934.3000 -6.3100 ;
        RECT 2799.0200 -9.3300 2802.0200 -6.3100 ;
        RECT -14.6800 104.1300 -11.6800 107.1500 ;
        RECT -14.6800 284.1300 -11.6800 287.1500 ;
        RECT -14.6800 464.1300 -11.6800 467.1500 ;
        RECT -14.6800 644.1300 -11.6800 647.1500 ;
        RECT -14.6800 824.1300 -11.6800 827.1500 ;
        RECT -14.6800 1004.1300 -11.6800 1007.1500 ;
        RECT -14.6800 1184.1300 -11.6800 1187.1500 ;
        RECT -14.6800 1364.1300 -11.6800 1367.1500 ;
        RECT -14.6800 1544.1300 -11.6800 1547.1500 ;
        RECT -14.6800 1724.1300 -11.6800 1727.1500 ;
        RECT 2931.3000 104.1300 2934.3000 107.1500 ;
        RECT 2931.3000 284.1300 2934.3000 287.1500 ;
        RECT 2931.3000 464.1300 2934.3000 467.1500 ;
        RECT 2931.3000 644.1300 2934.3000 647.1500 ;
        RECT 2931.3000 824.1300 2934.3000 827.1500 ;
        RECT 2931.3000 1004.1300 2934.3000 1007.1500 ;
        RECT 2931.3000 1184.1300 2934.3000 1187.1500 ;
        RECT 2931.3000 1364.1300 2934.3000 1367.1500 ;
        RECT 2931.3000 1544.1300 2934.3000 1547.1500 ;
        RECT 2931.3000 1724.1300 2934.3000 1727.1500 ;
        RECT -14.6800 1904.1300 -11.6800 1907.1500 ;
        RECT -14.6800 2084.1300 -11.6800 2087.1500 ;
        RECT -14.6800 2264.1300 -11.6800 2267.1500 ;
        RECT -14.6800 2444.1300 -11.6800 2447.1500 ;
        RECT -14.6800 2624.1300 -11.6800 2627.1500 ;
        RECT -14.6800 2804.1300 -11.6800 2807.1500 ;
        RECT -14.6800 2984.1300 -11.6800 2987.1500 ;
        RECT -14.6800 3164.1300 -11.6800 3167.1500 ;
        RECT -14.6800 3344.1300 -11.6800 3347.1500 ;
        RECT 2931.3000 1904.1300 2934.3000 1907.1500 ;
        RECT 2931.3000 2084.1300 2934.3000 2087.1500 ;
        RECT 2931.3000 2264.1300 2934.3000 2267.1500 ;
        RECT 2931.3000 2444.1300 2934.3000 2447.1500 ;
        RECT 2931.3000 2624.1300 2934.3000 2627.1500 ;
        RECT 2931.3000 2804.1300 2934.3000 2807.1500 ;
        RECT 2931.3000 2984.1300 2934.3000 2987.1500 ;
        RECT 2931.3000 3164.1300 2934.3000 3167.1500 ;
        RECT 2931.3000 3344.1300 2934.3000 3347.1500 ;
        RECT 99.0200 3525.9900 102.0200 3529.0100 ;
        RECT -14.6800 3525.9900 -11.6800 3529.0100 ;
        RECT 459.0200 3525.9900 462.0200 3529.0100 ;
        RECT 279.0200 3525.9900 282.0200 3529.0100 ;
        RECT 999.0200 3525.9900 1002.0200 3529.0100 ;
        RECT 819.0200 3525.9900 822.0200 3529.0100 ;
        RECT 639.0200 3525.9900 642.0200 3529.0100 ;
        RECT 1359.0200 3525.9900 1362.0200 3529.0100 ;
        RECT 1179.0200 3525.9900 1182.0200 3529.0100 ;
        RECT 1899.0200 3525.9900 1902.0200 3529.0100 ;
        RECT 1719.0200 3525.9900 1722.0200 3529.0100 ;
        RECT 1539.0200 3525.9900 1542.0200 3529.0100 ;
        RECT 2259.0200 3525.9900 2262.0200 3529.0100 ;
        RECT 2079.0200 3525.9900 2082.0200 3529.0100 ;
        RECT 2619.0200 3525.9900 2622.0200 3529.0100 ;
        RECT 2439.0200 3525.9900 2442.0200 3529.0100 ;
        RECT 2931.3000 3525.9900 2934.3000 3529.0100 ;
        RECT 2799.0200 3525.9900 2802.0200 3529.0100 ;
    END
# end of P/G power stripe data as pin

  END vssd1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 2917.6000 68.3800 2962.5000 71.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 68.3800 2.4000 71.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 248.3800 2962.5000 251.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 248.3800 2.4000 251.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 428.3800 2962.5000 431.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 428.3800 2.4000 431.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 608.3800 2962.5000 611.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 608.3800 2.4000 611.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 788.3800 2962.5000 791.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 788.3800 2.4000 791.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 968.3800 2962.5000 971.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 968.3800 2.4000 971.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1148.3800 2962.5000 1151.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1148.3800 2.4000 1151.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1328.3800 2962.5000 1331.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1328.3800 2.4000 1331.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1508.3800 2962.5000 1511.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1508.3800 2.4000 1511.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1688.3800 2962.5000 1691.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1688.3800 2.4000 1691.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1868.3800 2962.5000 1871.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 1868.3800 2.4000 1871.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2048.3800 2962.5000 2051.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2048.3800 2.4000 2051.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2228.3800 2962.5000 2231.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2228.3800 2.4000 2231.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2408.3800 2962.5000 2411.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2408.3800 2.4000 2411.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2588.3800 2962.5000 2591.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2588.3800 2.4000 2591.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2768.3800 2962.5000 2771.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2768.3800 2.4000 2771.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2948.3800 2962.5000 2951.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 2948.3800 2.4000 2951.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3128.3800 2962.5000 3131.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 3128.3800 2.4000 3131.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3308.3800 2962.5000 3311.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 3308.3800 2.4000 3311.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3488.3800 2962.5000 3491.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -42.8800 3488.3800 2.4000 3491.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.1800 3549.5000 2957.8000 3552.5000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2957.8000 -32.8200 2957.8000 -29.8200 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.0200 -37.5200 66.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.0200 3517.6000 66.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 243.0200 -37.5200 246.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 243.0200 3517.6000 246.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 423.0200 -37.5200 426.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 423.0200 3517.6000 426.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 603.0200 -37.5200 606.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 603.0200 3517.6000 606.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 783.0200 -37.5200 786.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 783.0200 3517.6000 786.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 963.0200 -37.5200 966.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 963.0200 3517.6000 966.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1143.0200 -37.5200 1146.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1143.0200 3517.6000 1146.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1323.0200 -37.5200 1326.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1323.0200 3517.6000 1326.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1503.0200 -37.5200 1506.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1503.0200 3517.6000 1506.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1683.0200 -37.5200 1686.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1683.0200 3517.6000 1686.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1863.0200 -37.5200 1866.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1863.0200 3517.6000 1866.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2043.0200 -37.5200 2046.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2043.0200 3517.6000 2046.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2223.0200 -37.5200 2226.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2223.0200 3517.6000 2226.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.0200 -37.5200 2406.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.0200 3517.6000 2406.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2583.0200 -37.5200 2586.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2583.0200 3517.6000 2586.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2763.0200 -37.5200 2766.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2763.0200 3517.6000 2766.0200 3557.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT -38.1800 3552.5000 -35.1800 3552.5000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2954.8000 -32.8200 2957.8000 3552.5000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT 2954.8000 -32.8200 2957.8000 3552.5000 ;
        RECT -38.1800 -32.8200 -35.1800 3552.5000 ;
      LAYER met5 ;
        RECT -38.1800 -32.8200 2957.8000 -29.8200 ;
        RECT -38.1800 3549.5000 2957.8000 3552.5000 ;
        RECT 63.0200 -32.8300 66.0200 -29.8100 ;
        RECT -38.1800 -32.8300 -35.1800 -29.8100 ;
        RECT 423.0200 -32.8300 426.0200 -29.8100 ;
        RECT 243.0200 -32.8300 246.0200 -29.8100 ;
        RECT 963.0200 -32.8300 966.0200 -29.8100 ;
        RECT 783.0200 -32.8300 786.0200 -29.8100 ;
        RECT 603.0200 -32.8300 606.0200 -29.8100 ;
        RECT 1323.0200 -32.8300 1326.0200 -29.8100 ;
        RECT 1143.0200 -32.8300 1146.0200 -29.8100 ;
        RECT 1863.0200 -32.8300 1866.0200 -29.8100 ;
        RECT 1683.0200 -32.8300 1686.0200 -29.8100 ;
        RECT 1503.0200 -32.8300 1506.0200 -29.8100 ;
        RECT 2223.0200 -32.8300 2226.0200 -29.8100 ;
        RECT 2043.0200 -32.8300 2046.0200 -29.8100 ;
        RECT 2583.0200 -32.8300 2586.0200 -29.8100 ;
        RECT 2763.0200 -32.8300 2766.0200 -29.8100 ;
        RECT 2403.0200 -32.8300 2406.0200 -29.8100 ;
        RECT 2954.8000 -32.8300 2957.8000 -29.8100 ;
        RECT -38.1800 68.3700 -35.1800 71.3900 ;
        RECT -38.1800 248.3700 -35.1800 251.3900 ;
        RECT -38.1800 428.3700 -35.1800 431.3900 ;
        RECT -38.1800 608.3700 -35.1800 611.3900 ;
        RECT -38.1800 788.3700 -35.1800 791.3900 ;
        RECT -38.1800 968.3700 -35.1800 971.3900 ;
        RECT -38.1800 1148.3700 -35.1800 1151.3900 ;
        RECT -38.1800 1328.3700 -35.1800 1331.3900 ;
        RECT -38.1800 1508.3700 -35.1800 1511.3900 ;
        RECT -38.1800 1688.3700 -35.1800 1691.3900 ;
        RECT 2954.8000 68.3700 2957.8000 71.3900 ;
        RECT 2954.8000 248.3700 2957.8000 251.3900 ;
        RECT 2954.8000 428.3700 2957.8000 431.3900 ;
        RECT 2954.8000 608.3700 2957.8000 611.3900 ;
        RECT 2954.8000 788.3700 2957.8000 791.3900 ;
        RECT 2954.8000 968.3700 2957.8000 971.3900 ;
        RECT 2954.8000 1148.3700 2957.8000 1151.3900 ;
        RECT 2954.8000 1328.3700 2957.8000 1331.3900 ;
        RECT 2954.8000 1508.3700 2957.8000 1511.3900 ;
        RECT 2954.8000 1688.3700 2957.8000 1691.3900 ;
        RECT -38.1800 1868.3700 -35.1800 1871.3900 ;
        RECT -38.1800 2048.3700 -35.1800 2051.3900 ;
        RECT -38.1800 2228.3700 -35.1800 2231.3900 ;
        RECT -38.1800 2408.3700 -35.1800 2411.3900 ;
        RECT -38.1800 2588.3700 -35.1800 2591.3900 ;
        RECT -38.1800 2768.3700 -35.1800 2771.3900 ;
        RECT -38.1800 2948.3700 -35.1800 2951.3900 ;
        RECT -38.1800 3128.3700 -35.1800 3131.3900 ;
        RECT -38.1800 3308.3700 -35.1800 3311.3900 ;
        RECT -38.1800 3488.3700 -35.1800 3491.3900 ;
        RECT 2954.8000 1868.3700 2957.8000 1871.3900 ;
        RECT 2954.8000 2048.3700 2957.8000 2051.3900 ;
        RECT 2954.8000 2228.3700 2957.8000 2231.3900 ;
        RECT 2954.8000 2408.3700 2957.8000 2411.3900 ;
        RECT 2954.8000 2588.3700 2957.8000 2591.3900 ;
        RECT 2954.8000 2768.3700 2957.8000 2771.3900 ;
        RECT 2954.8000 2948.3700 2957.8000 2951.3900 ;
        RECT 2954.8000 3128.3700 2957.8000 3131.3900 ;
        RECT 2954.8000 3308.3700 2957.8000 3311.3900 ;
        RECT 2954.8000 3488.3700 2957.8000 3491.3900 ;
        RECT 63.0200 3549.4900 66.0200 3552.5100 ;
        RECT -38.1800 3549.4900 -35.1800 3552.5100 ;
        RECT 423.0200 3549.4900 426.0200 3552.5100 ;
        RECT 243.0200 3549.4900 246.0200 3552.5100 ;
        RECT 963.0200 3549.4900 966.0200 3552.5100 ;
        RECT 783.0200 3549.4900 786.0200 3552.5100 ;
        RECT 603.0200 3549.4900 606.0200 3552.5100 ;
        RECT 1323.0200 3549.4900 1326.0200 3552.5100 ;
        RECT 1143.0200 3549.4900 1146.0200 3552.5100 ;
        RECT 1863.0200 3549.4900 1866.0200 3552.5100 ;
        RECT 1683.0200 3549.4900 1686.0200 3552.5100 ;
        RECT 1503.0200 3549.4900 1506.0200 3552.5100 ;
        RECT 2223.0200 3549.4900 2226.0200 3552.5100 ;
        RECT 2043.0200 3549.4900 2046.0200 3552.5100 ;
        RECT 2583.0200 3549.4900 2586.0200 3552.5100 ;
        RECT 2763.0200 3549.4900 2766.0200 3552.5100 ;
        RECT 2403.0200 3549.4900 2406.0200 3552.5100 ;
        RECT 2954.8000 3549.4900 2957.8000 3552.5100 ;
    END
# end of P/G power stripe data as pin

  END vdda2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 2917.6000 50.3800 2953.1000 53.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 50.3800 2.4000 53.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 230.3800 2953.1000 233.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 230.3800 2.4000 233.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 410.3800 2953.1000 413.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 410.3800 2.4000 413.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 590.3800 2953.1000 593.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 590.3800 2.4000 593.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 770.3800 2953.1000 773.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 770.3800 2.4000 773.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 950.3800 2953.1000 953.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 950.3800 2.4000 953.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1130.3800 2953.1000 1133.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1130.3800 2.4000 1133.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1310.3800 2953.1000 1313.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1310.3800 2.4000 1313.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1490.3800 2953.1000 1493.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1490.3800 2.4000 1493.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1670.3800 2953.1000 1673.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1670.3800 2.4000 1673.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1850.3800 2953.1000 1853.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 1850.3800 2.4000 1853.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2030.3800 2953.1000 2033.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2030.3800 2.4000 2033.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2210.3800 2953.1000 2213.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2210.3800 2.4000 2213.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2390.3800 2953.1000 2393.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2390.3800 2.4000 2393.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2570.3800 2953.1000 2573.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2570.3800 2.4000 2573.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2750.3800 2953.1000 2753.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2750.3800 2.4000 2753.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2930.3800 2953.1000 2933.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 2930.3800 2.4000 2933.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3110.3800 2953.1000 3113.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 3110.3800 2.4000 3113.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3290.3800 2953.1000 3293.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 3290.3800 2.4000 3293.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3470.3800 2953.1000 3473.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -33.4800 3470.3800 2.4000 3473.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -28.7800 3540.1000 2948.4000 3543.1000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2948.4000 -23.4200 2948.4000 -20.4200 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.0200 -28.1200 48.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.0200 3517.6000 48.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 225.0200 -28.1200 228.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 225.0200 3517.6000 228.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.0200 -28.1200 408.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.0200 3517.6000 408.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 585.0200 -28.1200 588.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 585.0200 3517.6000 588.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 765.0200 -28.1200 768.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 765.0200 3517.6000 768.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 945.0200 -28.1200 948.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 945.0200 3517.6000 948.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1125.0200 -28.1200 1128.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1125.0200 3517.6000 1128.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1305.0200 -28.1200 1308.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1305.0200 3517.6000 1308.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1485.0200 -28.1200 1488.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1485.0200 3517.6000 1488.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1665.0200 -28.1200 1668.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1665.0200 3517.6000 1668.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1845.0200 -28.1200 1848.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1845.0200 3517.6000 1848.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2025.0200 -28.1200 2028.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2025.0200 3517.6000 2028.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2205.0200 -28.1200 2208.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2205.0200 3517.6000 2208.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2385.0200 -28.1200 2388.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2385.0200 3517.6000 2388.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2565.0200 -28.1200 2568.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2565.0200 3517.6000 2568.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2745.0200 -28.1200 2748.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2745.0200 3517.6000 2748.0200 3547.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT -28.7800 3543.1000 -25.7800 3543.1000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2945.4000 -23.4200 2948.4000 3543.1000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT 2945.4000 -23.4200 2948.4000 3543.1000 ;
        RECT -28.7800 -23.4200 -25.7800 3543.1000 ;
      LAYER met5 ;
        RECT -28.7800 -23.4200 2948.4000 -20.4200 ;
        RECT -28.7800 3540.1000 2948.4000 3543.1000 ;
        RECT 45.0200 -23.4300 48.0200 -20.4100 ;
        RECT -28.7800 -23.4300 -25.7800 -20.4100 ;
        RECT 405.0200 -23.4300 408.0200 -20.4100 ;
        RECT 225.0200 -23.4300 228.0200 -20.4100 ;
        RECT 945.0200 -23.4300 948.0200 -20.4100 ;
        RECT 765.0200 -23.4300 768.0200 -20.4100 ;
        RECT 585.0200 -23.4300 588.0200 -20.4100 ;
        RECT 1305.0200 -23.4300 1308.0200 -20.4100 ;
        RECT 1125.0200 -23.4300 1128.0200 -20.4100 ;
        RECT 1845.0200 -23.4300 1848.0200 -20.4100 ;
        RECT 1665.0200 -23.4300 1668.0200 -20.4100 ;
        RECT 1485.0200 -23.4300 1488.0200 -20.4100 ;
        RECT 2205.0200 -23.4300 2208.0200 -20.4100 ;
        RECT 2025.0200 -23.4300 2028.0200 -20.4100 ;
        RECT 2745.0200 -23.4300 2748.0200 -20.4100 ;
        RECT 2565.0200 -23.4300 2568.0200 -20.4100 ;
        RECT 2385.0200 -23.4300 2388.0200 -20.4100 ;
        RECT 2945.4000 -23.4300 2948.4000 -20.4100 ;
        RECT -28.7800 50.3700 -25.7800 53.3900 ;
        RECT -28.7800 230.3700 -25.7800 233.3900 ;
        RECT -28.7800 410.3700 -25.7800 413.3900 ;
        RECT -28.7800 590.3700 -25.7800 593.3900 ;
        RECT -28.7800 770.3700 -25.7800 773.3900 ;
        RECT -28.7800 950.3700 -25.7800 953.3900 ;
        RECT -28.7800 1130.3700 -25.7800 1133.3900 ;
        RECT -28.7800 1310.3700 -25.7800 1313.3900 ;
        RECT -28.7800 1490.3700 -25.7800 1493.3900 ;
        RECT -28.7800 1670.3700 -25.7800 1673.3900 ;
        RECT 2945.4000 50.3700 2948.4000 53.3900 ;
        RECT 2945.4000 230.3700 2948.4000 233.3900 ;
        RECT 2945.4000 410.3700 2948.4000 413.3900 ;
        RECT 2945.4000 590.3700 2948.4000 593.3900 ;
        RECT 2945.4000 770.3700 2948.4000 773.3900 ;
        RECT 2945.4000 950.3700 2948.4000 953.3900 ;
        RECT 2945.4000 1130.3700 2948.4000 1133.3900 ;
        RECT 2945.4000 1310.3700 2948.4000 1313.3900 ;
        RECT 2945.4000 1490.3700 2948.4000 1493.3900 ;
        RECT 2945.4000 1670.3700 2948.4000 1673.3900 ;
        RECT -28.7800 1850.3700 -25.7800 1853.3900 ;
        RECT -28.7800 2030.3700 -25.7800 2033.3900 ;
        RECT -28.7800 2210.3700 -25.7800 2213.3900 ;
        RECT -28.7800 2390.3700 -25.7800 2393.3900 ;
        RECT -28.7800 2570.3700 -25.7800 2573.3900 ;
        RECT -28.7800 2750.3700 -25.7800 2753.3900 ;
        RECT -28.7800 2930.3700 -25.7800 2933.3900 ;
        RECT -28.7800 3110.3700 -25.7800 3113.3900 ;
        RECT -28.7800 3290.3700 -25.7800 3293.3900 ;
        RECT -28.7800 3470.3700 -25.7800 3473.3900 ;
        RECT 2945.4000 1850.3700 2948.4000 1853.3900 ;
        RECT 2945.4000 2030.3700 2948.4000 2033.3900 ;
        RECT 2945.4000 2210.3700 2948.4000 2213.3900 ;
        RECT 2945.4000 2390.3700 2948.4000 2393.3900 ;
        RECT 2945.4000 2570.3700 2948.4000 2573.3900 ;
        RECT 2945.4000 2750.3700 2948.4000 2753.3900 ;
        RECT 2945.4000 2930.3700 2948.4000 2933.3900 ;
        RECT 2945.4000 3110.3700 2948.4000 3113.3900 ;
        RECT 2945.4000 3290.3700 2948.4000 3293.3900 ;
        RECT 2945.4000 3470.3700 2948.4000 3473.3900 ;
        RECT 45.0200 3540.0900 48.0200 3543.1100 ;
        RECT -28.7800 3540.0900 -25.7800 3543.1100 ;
        RECT 405.0200 3540.0900 408.0200 3543.1100 ;
        RECT 225.0200 3540.0900 228.0200 3543.1100 ;
        RECT 945.0200 3540.0900 948.0200 3543.1100 ;
        RECT 765.0200 3540.0900 768.0200 3543.1100 ;
        RECT 585.0200 3540.0900 588.0200 3543.1100 ;
        RECT 1305.0200 3540.0900 1308.0200 3543.1100 ;
        RECT 1125.0200 3540.0900 1128.0200 3543.1100 ;
        RECT 1845.0200 3540.0900 1848.0200 3543.1100 ;
        RECT 1665.0200 3540.0900 1668.0200 3543.1100 ;
        RECT 1485.0200 3540.0900 1488.0200 3543.1100 ;
        RECT 2205.0200 3540.0900 2208.0200 3543.1100 ;
        RECT 2025.0200 3540.0900 2028.0200 3543.1100 ;
        RECT 2745.0200 3540.0900 2748.0200 3543.1100 ;
        RECT 2565.0200 3540.0900 2568.0200 3543.1100 ;
        RECT 2385.0200 3540.0900 2388.0200 3543.1100 ;
        RECT 2945.4000 3540.0900 2948.4000 3543.1100 ;
    END
# end of P/G power stripe data as pin

  END vdda1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 2917.6000 32.3800 2943.7000 35.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 32.3800 2.4000 35.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 212.3800 2943.7000 215.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 212.3800 2.4000 215.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 392.3800 2943.7000 395.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 392.3800 2.4000 395.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 572.3800 2943.7000 575.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 572.3800 2.4000 575.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 752.3800 2943.7000 755.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 752.3800 2.4000 755.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 932.3800 2943.7000 935.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 932.3800 2.4000 935.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1112.3800 2943.7000 1115.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1112.3800 2.4000 1115.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1292.3800 2943.7000 1295.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1292.3800 2.4000 1295.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1472.3800 2943.7000 1475.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1472.3800 2.4000 1475.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1652.3800 2943.7000 1655.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1652.3800 2.4000 1655.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1832.3800 2943.7000 1835.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 1832.3800 2.4000 1835.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2012.3800 2943.7000 2015.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2012.3800 2.4000 2015.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2192.3800 2943.7000 2195.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2192.3800 2.4000 2195.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2372.3800 2943.7000 2375.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2372.3800 2.4000 2375.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2552.3800 2943.7000 2555.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2552.3800 2.4000 2555.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2732.3800 2943.7000 2735.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2732.3800 2.4000 2735.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2912.3800 2943.7000 2915.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 2912.3800 2.4000 2915.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3092.3800 2943.7000 3095.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 3092.3800 2.4000 3095.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3272.3800 2943.7000 3275.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 3272.3800 2.4000 3275.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3452.3800 2943.7000 3455.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.0800 3452.3800 2.4000 3455.3800 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.3800 3530.7000 2939.0000 3533.7000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2939.0000 -14.0200 2939.0000 -11.0200 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.0200 -18.7200 30.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.0200 3517.6000 30.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 207.0200 -18.7200 210.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 207.0200 3517.6000 210.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.0200 -18.7200 390.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.0200 3517.6000 390.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.0200 -18.7200 570.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.0200 3517.6000 570.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 747.0200 -18.7200 750.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 747.0200 3517.6000 750.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.0200 -18.7200 930.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.0200 3517.6000 930.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.0200 -18.7200 1110.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.0200 3517.6000 1110.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.0200 -18.7200 1290.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.0200 3517.6000 1290.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1467.0200 -18.7200 1470.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1467.0200 3517.6000 1470.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1647.0200 -18.7200 1650.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1647.0200 3517.6000 1650.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.0200 -18.7200 1830.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.0200 3517.6000 1830.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.0200 -18.7200 2010.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.0200 3517.6000 2010.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.0200 -18.7200 2190.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.0200 3517.6000 2190.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2367.0200 -18.7200 2370.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2367.0200 3517.6000 2370.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.0200 -18.7200 2550.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.0200 3517.6000 2550.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2727.0200 -18.7200 2730.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2727.0200 3517.6000 2730.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2907.0200 -18.7200 2910.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2907.0200 3517.6000 2910.0200 3538.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT -19.3800 3533.7000 -16.3800 3533.7000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2936.0000 -14.0200 2939.0000 3533.7000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT 2936.0000 -14.0200 2939.0000 3533.7000 ;
        RECT -19.3800 -14.0200 -16.3800 3533.7000 ;
      LAYER met5 ;
        RECT -19.3800 -14.0200 2939.0000 -11.0200 ;
        RECT -19.3800 3530.7000 2939.0000 3533.7000 ;
        RECT 27.0200 -14.0300 30.0200 -11.0100 ;
        RECT -19.3800 -14.0300 -16.3800 -11.0100 ;
        RECT 567.0200 -14.0300 570.0200 -11.0100 ;
        RECT 387.0200 -14.0300 390.0200 -11.0100 ;
        RECT 207.0200 -14.0300 210.0200 -11.0100 ;
        RECT 747.0200 -14.0300 750.0200 -11.0100 ;
        RECT 927.0200 -14.0300 930.0200 -11.0100 ;
        RECT 1107.0200 -14.0300 1110.0200 -11.0100 ;
        RECT 1287.0200 -14.0300 1290.0200 -11.0100 ;
        RECT 1467.0200 -14.0300 1470.0200 -11.0100 ;
        RECT 1647.0200 -14.0300 1650.0200 -11.0100 ;
        RECT 1827.0200 -14.0300 1830.0200 -11.0100 ;
        RECT 2007.0200 -14.0300 2010.0200 -11.0100 ;
        RECT 2187.0200 -14.0300 2190.0200 -11.0100 ;
        RECT 2367.0200 -14.0300 2370.0200 -11.0100 ;
        RECT 2547.0200 -14.0300 2550.0200 -11.0100 ;
        RECT 2727.0200 -14.0300 2730.0200 -11.0100 ;
        RECT 2907.0200 -14.0300 2910.0200 -11.0100 ;
        RECT 2936.0000 -14.0300 2939.0000 -11.0100 ;
        RECT -19.3800 32.3700 -16.3800 35.3900 ;
        RECT -19.3800 212.3700 -16.3800 215.3900 ;
        RECT -19.3800 392.3700 -16.3800 395.3900 ;
        RECT -19.3800 572.3700 -16.3800 575.3900 ;
        RECT -19.3800 752.3700 -16.3800 755.3900 ;
        RECT -19.3800 932.3700 -16.3800 935.3900 ;
        RECT -19.3800 1112.3700 -16.3800 1115.3900 ;
        RECT -19.3800 1292.3700 -16.3800 1295.3900 ;
        RECT -19.3800 1472.3700 -16.3800 1475.3900 ;
        RECT -19.3800 1652.3700 -16.3800 1655.3900 ;
        RECT 2936.0000 32.3700 2939.0000 35.3900 ;
        RECT 2936.0000 212.3700 2939.0000 215.3900 ;
        RECT 2936.0000 392.3700 2939.0000 395.3900 ;
        RECT 2936.0000 572.3700 2939.0000 575.3900 ;
        RECT 2936.0000 752.3700 2939.0000 755.3900 ;
        RECT 2936.0000 932.3700 2939.0000 935.3900 ;
        RECT 2936.0000 1112.3700 2939.0000 1115.3900 ;
        RECT 2936.0000 1292.3700 2939.0000 1295.3900 ;
        RECT 2936.0000 1472.3700 2939.0000 1475.3900 ;
        RECT 2936.0000 1652.3700 2939.0000 1655.3900 ;
        RECT -19.3800 1832.3700 -16.3800 1835.3900 ;
        RECT -19.3800 2012.3700 -16.3800 2015.3900 ;
        RECT -19.3800 2192.3700 -16.3800 2195.3900 ;
        RECT -19.3800 2372.3700 -16.3800 2375.3900 ;
        RECT -19.3800 2552.3700 -16.3800 2555.3900 ;
        RECT -19.3800 2732.3700 -16.3800 2735.3900 ;
        RECT -19.3800 2912.3700 -16.3800 2915.3900 ;
        RECT -19.3800 3092.3700 -16.3800 3095.3900 ;
        RECT -19.3800 3272.3700 -16.3800 3275.3900 ;
        RECT -19.3800 3452.3700 -16.3800 3455.3900 ;
        RECT 2936.0000 1832.3700 2939.0000 1835.3900 ;
        RECT 2936.0000 2012.3700 2939.0000 2015.3900 ;
        RECT 2936.0000 2192.3700 2939.0000 2195.3900 ;
        RECT 2936.0000 2372.3700 2939.0000 2375.3900 ;
        RECT 2936.0000 2552.3700 2939.0000 2555.3900 ;
        RECT 2936.0000 2732.3700 2939.0000 2735.3900 ;
        RECT 2936.0000 2912.3700 2939.0000 2915.3900 ;
        RECT 2936.0000 3092.3700 2939.0000 3095.3900 ;
        RECT 2936.0000 3272.3700 2939.0000 3275.3900 ;
        RECT 2936.0000 3452.3700 2939.0000 3455.3900 ;
        RECT 27.0200 3530.6900 30.0200 3533.7100 ;
        RECT -19.3800 3530.6900 -16.3800 3533.7100 ;
        RECT 567.0200 3530.6900 570.0200 3533.7100 ;
        RECT 387.0200 3530.6900 390.0200 3533.7100 ;
        RECT 207.0200 3530.6900 210.0200 3533.7100 ;
        RECT 927.0200 3530.6900 930.0200 3533.7100 ;
        RECT 747.0200 3530.6900 750.0200 3533.7100 ;
        RECT 1107.0200 3530.6900 1110.0200 3533.7100 ;
        RECT 1287.0200 3530.6900 1290.0200 3533.7100 ;
        RECT 1467.0200 3530.6900 1470.0200 3533.7100 ;
        RECT 1647.0200 3530.6900 1650.0200 3533.7100 ;
        RECT 1827.0200 3530.6900 1830.0200 3533.7100 ;
        RECT 2007.0200 3530.6900 2010.0200 3533.7100 ;
        RECT 2187.0200 3530.6900 2190.0200 3533.7100 ;
        RECT 2367.0200 3530.6900 2370.0200 3533.7100 ;
        RECT 2547.0200 3530.6900 2550.0200 3533.7100 ;
        RECT 2727.0200 3530.6900 2730.0200 3533.7100 ;
        RECT 2907.0200 3530.6900 2910.0200 3533.7100 ;
        RECT 2936.0000 3530.6900 2939.0000 3533.7100 ;
    END
# end of P/G power stripe data as pin

  END vccd2
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 2917.6000 14.1400 2934.3000 17.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 14.1400 2.4000 17.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 194.1400 2934.3000 197.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 194.1400 2.4000 197.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 374.1400 2934.3000 377.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 374.1400 2.4000 377.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 554.1400 2934.3000 557.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 554.1400 2.4000 557.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 734.1400 2934.3000 737.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 734.1400 2.4000 737.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 914.1400 2934.3000 917.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 914.1400 2.4000 917.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1094.1400 2934.3000 1097.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1094.1400 2.4000 1097.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1274.1400 2934.3000 1277.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1274.1400 2.4000 1277.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1454.1400 2934.3000 1457.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1454.1400 2.4000 1457.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1634.1400 2934.3000 1637.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1634.1400 2.4000 1637.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1814.1400 2934.3000 1817.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1814.1400 2.4000 1817.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 1994.1400 2934.3000 1997.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 1994.1400 2.4000 1997.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2174.1400 2934.3000 2177.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2174.1400 2.4000 2177.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2354.1400 2934.3000 2357.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2354.1400 2.4000 2357.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2534.1400 2934.3000 2537.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2534.1400 2.4000 2537.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2714.1400 2934.3000 2717.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2714.1400 2.4000 2717.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 2894.1400 2934.3000 2897.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 2894.1400 2.4000 2897.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3074.1400 2934.3000 3077.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 3074.1400 2.4000 3077.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3254.1400 2934.3000 3257.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 3254.1400 2.4000 3257.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT 2917.6000 3434.1400 2934.3000 3437.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.6800 3434.1400 2.4000 3437.1400 ;
    END
    PORT
      LAYER met5 ;
        RECT -9.9800 3521.3000 2929.6000 3524.3000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2929.6000 -4.6200 2929.6000 -1.6200 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.0200 -9.3200 12.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.0200 3517.6000 12.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 189.0200 -9.3200 192.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 189.0200 3517.6000 192.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 369.0200 -9.3200 372.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 369.0200 3517.6000 372.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 549.0200 -9.3200 552.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 549.0200 3517.6000 552.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 729.0200 -9.3200 732.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 729.0200 3517.6000 732.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 909.0200 -9.3200 912.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 909.0200 3517.6000 912.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1089.0200 -9.3200 1092.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1089.0200 3517.6000 1092.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1269.0200 -9.3200 1272.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1269.0200 3517.6000 1272.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1449.0200 -9.3200 1452.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1449.0200 3517.6000 1452.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1629.0200 -9.3200 1632.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1629.0200 3517.6000 1632.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1809.0200 -9.3200 1812.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1809.0200 3517.6000 1812.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1989.0200 -9.3200 1992.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1989.0200 3517.6000 1992.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2169.0200 -9.3200 2172.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2169.0200 3517.6000 2172.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2349.0200 -9.3200 2352.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2349.0200 3517.6000 2352.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2529.0200 -9.3200 2532.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2529.0200 3517.6000 2532.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.0200 -9.3200 2712.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.0200 3517.6000 2712.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2889.0200 -9.3200 2892.0200 2.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2889.0200 3517.6000 2892.0200 3529.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT -9.9800 3524.3000 -6.9800 3524.3000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2926.6000 -4.6200 2929.6000 3524.3000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT 2926.6000 -4.6200 2929.6000 3524.3000 ;
        RECT -9.9800 -4.6200 -6.9800 3524.3000 ;
        RECT 549.0200 0.0000 552.0200 3520.0000 ;
        RECT 369.0200 0.0000 372.0200 3520.0000 ;
        RECT 189.0200 0.0000 192.0200 3520.0000 ;
        RECT 9.0200 0.0000 12.0200 3520.0000 ;
        RECT 1449.0200 0.0000 1452.0200 3520.0000 ;
        RECT 1269.0200 0.0000 1272.0200 3520.0000 ;
        RECT 1089.0200 0.0000 1092.0200 3520.0000 ;
        RECT 909.0200 0.0000 912.0200 3520.0000 ;
        RECT 729.0200 0.0000 732.0200 3520.0000 ;
        RECT 2169.0200 0.0000 2172.0200 3520.0000 ;
        RECT 1989.0200 0.0000 1992.0200 3520.0000 ;
        RECT 1809.0200 0.0000 1812.0200 3520.0000 ;
        RECT 1629.0200 0.0000 1632.0200 3520.0000 ;
        RECT 2889.0200 0.0000 2892.0200 3520.0000 ;
        RECT 2709.0200 0.0000 2712.0200 3520.0000 ;
        RECT 2529.0200 0.0000 2532.0200 3520.0000 ;
        RECT 2349.0200 0.0000 2352.0200 3520.0000 ;
      LAYER met5 ;
        RECT -9.9800 -4.6200 2929.6000 -1.6200 ;
        RECT 0.0000 14.1400 2920.0000 17.1400 ;
        RECT 0.0000 194.1400 2920.0000 197.1400 ;
        RECT 0.0000 374.1400 2920.0000 377.1400 ;
        RECT 0.0000 554.1400 2920.0000 557.1400 ;
        RECT 0.0000 734.1400 2920.0000 737.1400 ;
        RECT 0.0000 914.1400 2920.0000 917.1400 ;
        RECT 0.0000 1094.1400 2920.0000 1097.1400 ;
        RECT 0.0000 1274.1400 2920.0000 1277.1400 ;
        RECT 0.0000 1454.1400 2920.0000 1457.1400 ;
        RECT 0.0000 1634.1400 2920.0000 1637.1400 ;
        RECT 0.0000 1814.1400 2920.0000 1817.1400 ;
        RECT 0.0000 1994.1400 2920.0000 1997.1400 ;
        RECT 0.0000 2174.1400 2920.0000 2177.1400 ;
        RECT 0.0000 2354.1400 2920.0000 2357.1400 ;
        RECT 0.0000 2534.1400 2920.0000 2537.1400 ;
        RECT 0.0000 2714.1400 2920.0000 2717.1400 ;
        RECT 0.0000 2894.1400 2920.0000 2897.1400 ;
        RECT 0.0000 3074.1400 2920.0000 3077.1400 ;
        RECT 0.0000 3254.1400 2920.0000 3257.1400 ;
        RECT 0.0000 3434.1400 2920.0000 3437.1400 ;
        RECT -9.9800 3521.3000 2929.6000 3524.3000 ;
        RECT -9.9800 -4.6300 -6.9800 -1.6100 ;
        RECT 9.0200 -4.6300 12.0200 -1.6100 ;
        RECT 189.0200 -4.6300 192.0200 -1.6100 ;
        RECT 369.0200 -4.6300 372.0200 -1.6100 ;
        RECT 549.0200 -4.6300 552.0200 -1.6100 ;
        RECT 729.0200 -4.6300 732.0200 -1.6100 ;
        RECT 909.0200 -4.6300 912.0200 -1.6100 ;
        RECT 1089.0200 -4.6300 1092.0200 -1.6100 ;
        RECT 1269.0200 -4.6300 1272.0200 -1.6100 ;
        RECT 1449.0200 -4.6300 1452.0200 -1.6100 ;
        RECT 1629.0200 -4.6300 1632.0200 -1.6100 ;
        RECT 1809.0200 -4.6300 1812.0200 -1.6100 ;
        RECT 1989.0200 -4.6300 1992.0200 -1.6100 ;
        RECT 2169.0200 -4.6300 2172.0200 -1.6100 ;
        RECT 2349.0200 -4.6300 2352.0200 -1.6100 ;
        RECT 2529.0200 -4.6300 2532.0200 -1.6100 ;
        RECT 2709.0200 -4.6300 2712.0200 -1.6100 ;
        RECT 2889.0200 -4.6300 2892.0200 -1.6100 ;
        RECT 2926.6000 -4.6300 2929.6000 -1.6100 ;
        RECT -9.9800 14.1300 -6.9800 17.1500 ;
        RECT -9.9800 194.1300 -6.9800 197.1500 ;
        RECT -9.9800 374.1300 -6.9800 377.1500 ;
        RECT -9.9800 554.1300 -6.9800 557.1500 ;
        RECT -9.9800 734.1300 -6.9800 737.1500 ;
        RECT -9.9800 914.1300 -6.9800 917.1500 ;
        RECT -9.9800 1094.1300 -6.9800 1097.1500 ;
        RECT -9.9800 1274.1300 -6.9800 1277.1500 ;
        RECT -9.9800 1454.1300 -6.9800 1457.1500 ;
        RECT -9.9800 1634.1300 -6.9800 1637.1500 ;
        RECT 2926.6000 14.1300 2929.6000 17.1500 ;
        RECT 2926.6000 194.1300 2929.6000 197.1500 ;
        RECT 2926.6000 374.1300 2929.6000 377.1500 ;
        RECT 2926.6000 554.1300 2929.6000 557.1500 ;
        RECT 2926.6000 734.1300 2929.6000 737.1500 ;
        RECT 2926.6000 914.1300 2929.6000 917.1500 ;
        RECT 2926.6000 1094.1300 2929.6000 1097.1500 ;
        RECT 2926.6000 1274.1300 2929.6000 1277.1500 ;
        RECT 2926.6000 1454.1300 2929.6000 1457.1500 ;
        RECT 2926.6000 1634.1300 2929.6000 1637.1500 ;
        RECT -9.9800 1814.1300 -6.9800 1817.1500 ;
        RECT -9.9800 1994.1300 -6.9800 1997.1500 ;
        RECT -9.9800 2174.1300 -6.9800 2177.1500 ;
        RECT -9.9800 2354.1300 -6.9800 2357.1500 ;
        RECT -9.9800 2534.1300 -6.9800 2537.1500 ;
        RECT -9.9800 2714.1300 -6.9800 2717.1500 ;
        RECT -9.9800 2894.1300 -6.9800 2897.1500 ;
        RECT -9.9800 3074.1300 -6.9800 3077.1500 ;
        RECT -9.9800 3254.1300 -6.9800 3257.1500 ;
        RECT -9.9800 3434.1300 -6.9800 3437.1500 ;
        RECT 2926.6000 1814.1300 2929.6000 1817.1500 ;
        RECT 2926.6000 1994.1300 2929.6000 1997.1500 ;
        RECT 2926.6000 2174.1300 2929.6000 2177.1500 ;
        RECT 2926.6000 2354.1300 2929.6000 2357.1500 ;
        RECT 2926.6000 2534.1300 2929.6000 2537.1500 ;
        RECT 2926.6000 2714.1300 2929.6000 2717.1500 ;
        RECT 2926.6000 2894.1300 2929.6000 2897.1500 ;
        RECT 2926.6000 3074.1300 2929.6000 3077.1500 ;
        RECT 2926.6000 3254.1300 2929.6000 3257.1500 ;
        RECT 2926.6000 3434.1300 2929.6000 3437.1500 ;
        RECT -9.9800 3521.2900 -6.9800 3524.3100 ;
        RECT 9.0200 3521.2900 12.0200 3524.3100 ;
        RECT 189.0200 3521.2900 192.0200 3524.3100 ;
        RECT 369.0200 3521.2900 372.0200 3524.3100 ;
        RECT 549.0200 3521.2900 552.0200 3524.3100 ;
        RECT 729.0200 3521.2900 732.0200 3524.3100 ;
        RECT 909.0200 3521.2900 912.0200 3524.3100 ;
        RECT 1089.0200 3521.2900 1092.0200 3524.3100 ;
        RECT 1269.0200 3521.2900 1272.0200 3524.3100 ;
        RECT 1449.0200 3521.2900 1452.0200 3524.3100 ;
        RECT 1629.0200 3521.2900 1632.0200 3524.3100 ;
        RECT 1809.0200 3521.2900 1812.0200 3524.3100 ;
        RECT 1989.0200 3521.2900 1992.0200 3524.3100 ;
        RECT 2169.0200 3521.2900 2172.0200 3524.3100 ;
        RECT 2349.0200 3521.2900 2352.0200 3524.3100 ;
        RECT 2529.0200 3521.2900 2532.0200 3524.3100 ;
        RECT 2709.0200 3521.2900 2712.0200 3524.3100 ;
        RECT 2889.0200 3521.2900 2892.0200 3524.3100 ;
        RECT 2926.6000 3521.2900 2929.6000 3524.3100 ;
    END
# end of P/G power stripe data as pin

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.0000 0.0000 2920.0000 3520.0000 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 2920.0000 3520.0000 ;
    LAYER met2 ;
      RECT 0.0000 0.0000 2920.0000 3520.0000 ;
    LAYER met3 ;
      RECT 0.0000 0.0000 2920.0000 3520.0000 ;
    LAYER met4 ;
      RECT 0.0000 0.0000 2920.0000 3520.0000 ;
    LAYER met5 ;
      RECT 0.0000 0.0000 2920.0000 3520.0000 ;
  END
END user_project_wrapper

END LIBRARY
